                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����tJ xS[   	��!$�	 �:   %��!�9D ��   ���!��� �W U��{�
ˇX�0�4�5�G�  ���������������������������������� ��  ���� �$  
� ��  �� �   
� ��  ��  � 0�  
� ��  �� �   
  � ��  ��  � 0�  
� ��  �� �   
  � �� @�� �� P��`�� T��| ��  ��  � 0�     �h ��h��h0�� P�  
 Q� �4 �4���:P��  �� S� �4���:  ����� � � �����  $ ���D*D*D*D*p@-�1  �p@��4  ��P � � `�� ���  �  U�  6  �  P�  x ��x��	�� � �����l ��d��	������  �  V�  
T ��H��	������  �_ � P�  8 ��(��	������  �( ����	�� � �����  ��p���` ��  �P�P�P�P�P�Pa �ި ��	��p�� ���/� �����  
 ���/�  ������ � �����0@-� 0��h ���G��  ��  �\ ����  Q�     �QX��!��QT�� ���P� �� 0�� � � ��� �  R����: T�  
  ��0��� ������   � P@-� @��`����< �� ��2�/� P�   �����  ������@-� @��,����D �� ��2�/� P�   �����  ������@-����l ��0�/����p@-� @��������T�����*����00�� ��3�/� P�   ��p���  ������@-����� @����*����X0�� ��3�/�  P�  
 �����  ������@-�h��p ��0�/����@-�T����` ��
��2�/� �����@-����� @��,��*����d0�� ��3�/�  P�  
��h ��0�/�  P�  
 �����  ������  �������C-� @��  ��  �� P����� ���i�����P�� ��1�/� �� ��^ � P�� �� ��Z � p�� � �	  � �� �����%
��t��L0�� ��3�/�@�� T����: ������@-� @�� T�B  
  � T��0�  �C  �8  �.  �8  �A  �L  �@  �+  �W  �]  �N  �h  �z  �y  �r  �w  �7  �+  � T�G  

  � D� P� �0n  �%  �.  �8  �-  �  �C  �I  � T�+  
  � T�Q  
 T�$  
 T�^  "  �T�O  
�� ��  
 P�V  <  � � � � � � � � �Y���  P�   ���O  � � � � � � � � � � �0���  P�   ���E  � � � � � � � � � � � � � � � � � � �/���  P�   ����7  � � � � �}���  P�   ����0  � � � � �D���  P�   ����)  � � � � �  �  P�   ����"  � � � � �  �  P�   ����  � � �D���  P�   ����  � � � � �E���  P�   ����  � � �2���  P�   ����  � � ����  P�   ����  � � ����� � � � � �����  �@-����� `��T��!Z��<�� 0��(0��+��C� ��  � @��  T�   ������  ������ ��G-� @��P��`��p��(���3�����0�� ��C�� ��0���<�/� ���  Y�  
	 ������  �������@-�t�� ���l����� �`����0�T����@�H����P�<����`�0�����p�(������  Q�B  
  R�   ��?  � S�   T�   T�    W�    \�   ��3  � ��1  �  W�   \�   ��+  � ��)  �  U�    V�   T�    W�    \�   ��  � ��  �  W�   \�   ��  � ��  � T�    W�    \�   ��  � ��	  �  W�   \�   � � � ����� ��   �  ������     p@-�P�� @��  ��� �� � P�   ��p���@�� T�����  ������p@-�P�� @��  ��� �� � P�   ��p���@�� T�����  �������O-�  ��
���@���P���`���p����������؀��ܐ����� �� ��T
��� �� ��H
��� ��  �� 0��  ���4 ���� ��0�� S����: 0��  ���5 ���� ��0�� S����: 0��  ���6 ���� ��0�� S����: 0��  ���7 ���� ��0�� S����: 0��  ���< ���� ��0�� S����: 0��  ���> ���� ��0�� S����: 0��  ���8 ���� ��0�� S����: 0��  ���9 ���� ��0�� S����: 0��  ���: ���  � ��0�� S����: 0��  ������; ���  � ��0�� S����: 0��  ������; ���  � ��0�� S����: 0��  ��� ���; ���  � ��0�� S����: �������C-��M� @��P��h��@ ���p �  W�   ��ݍ����� W�  �  ������ U�  
 U�    � � �������  � � �������  � � �  ������ � ���� ��V���  P�    ������ `��  �� ����	�� P�  *� ����  ����  ������ ��  �  ������`�� V����: ������|��  ����  ���/�h��  ����  ���/�T��  ����  ���/�  ��'����4'��P���/�@-�p ���F�� �� 0��   �0�� �  S����:p ���F�� �� ��	  ���� ��@ �  
  ���F�� �� ����������  Q����:  ������ ��  ����( �� �  
 ���/�����  Q����:  �������O-� @��P��`��p��  �� �婉� V�  
 V�    � � ���������  �����	  � � ���������  �����  � � �  ������ � �  �����( ����� �� �� ������� W�  � ��   � �� �� ����� �� ��( �������0 ����� �� ����� �� ��( ��  �� �� ��  �  ����� �� �� �� �� ��	 P����:  �� ��  � ����5 ���  ���� �� �� �� �� ��
 P����: V�  
0 ����� ��  W�  ����  P�  ����� W�  � ��   � �� �� ����� ��  �����b���  P�  ����� W�  � ��   � �� �� ����� ��  ����� �����( ����� �� �� ����� ��0 �� ����  �� ����  �� V�  
 ��9���3���-���  �� ��  ���� �� �� �� �� �� �� �� P����:  �� ��  ���� �� �� �� �� �� P����: V�   
������ �� ����� �� � ���0 ������
����0 �� � �|��0 ������ �� D������  P�  ����� W�  � ��   � �� �� ����� ��  ��F������( ��  �  
  �����( ������� W�  � ��   � �� �� ����� ��  ��2�������� W�  � ��   � �� �� ����� �� ��%����O-� @��P��`��p�������  ����x��  �� W�   ��  �� �� ��  ����� W�  H��  �� �� ��8��  �����,��  ����J�����  ��
�� ���  � ���
�� A�
���  �  �����
  � ��	�� ��(0������  P�    ������
������  �� ��	 P����� ������@-� @������� T�  � ��   � �� �� ����� �� ��( ��  �� ��� �� ��  T�  ����  P�  ����� T�  � ��   � �� �� ����� ��  �����w���  P�  ����� T�  � ��   � �� �� ����� ��  ����������� T�  � ��   � �� �� ����� �� ������@-� @��r����  �� �� �� �����  P�    ����� �������C-� @��P��X`����� ���y�� ������  P�    ������0�� ���� �� P��\���  P�    ������ ������  � Zb P0��!  J  ��0q�  : 2q�  : 4q�  : ���   �3q��@  �� 3q�@  ��2q��@  �� 2q�@  ��1q��@  �� 1q�@  ��0q�� @  ��P� �1 ���/�!� aB@�2�  `" 2q�  : 4q�  :�� 4q�?#��  :�� 4q�?&��  :�� 4q�?)���!?,�# 0q�  *!�!�3q��@  �� 3q�@  ��2q��@  �� 2q�@  ��1q��@  �� 1q�@  �����*�0q�� @  ��P� �1 ���ϰ�  `B a"�/��ϰ�  `B@-�  ��  �����  �� 2q���: 4q���: �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    20120823                                                a  � � �L5l5D    � � � �	  �����y  ���������������������D    4$ş� �0� ���!�1 ��/�՟��o��� � � � � � � � � � � � � � � � ��V �` �%h�� V��������  6�! 6" 60�@��0�0 V�0�����0��0�����0����Q�����Q�0� ��0���l��T����T����0�A ��0���L����� �� $�� ��������!���������������!� ��  ����������������������� ��� �������!�  �����
�� �� �������!������  ��������������!���� ��� ��#�� Q�  
�  �  ��� �x  ����}  �  �t  ����� p�  
� p�   
� p�6  
� p�N  
R   @-� Q�	  
  Q�
  
 Q�  
 Q�  
@ Q�  
 @��G  � � @��D  � � @��A  �. � @��>  �B � @��;  �] � @��8  ���1����6  ����/�� ��������������(����� Q�D � �����!�����  ����p��0����/�� ��,  �  P�  
X���� ������d��������������(��� �����!�d �� ��� ���� @-�5 � @��  �����  ����  ���� @-� Q��    Q�   Q��   Q��  @ Q�  @����        ������!��':��  ���� �� ������������!��1������8!��01������8!��01������8!��01��x����8!��01����H���� �����������L��������(��<��������(��,��������(����������(����������(�����(����,����� ���� �������� �� ������������� ���� ������� �� ���� ���� ������� �� ���� ���� ������� �� ������ P �  P   �$���   �    � p��  p  q  r  s            H  I @H @I �H �I �H �I � � � � � � H-�����M� �0�0��  S�  
0�0�� ��0� 0����0� ��0�0��0c� ��0� ���0�0�����0�0��0c�̠� ���# � 0��  S�   
�����K� ��� H-���� �M� ��  �  �0K� �� �� ��00 �2@� 0�� �� �3�/�  ������K� ��� H-���� �M� ��  �  �0K� �� �� ��40 �2@� 0�� �� �3�/�  �����K� ��� H-�����M� �� � �0K� �� �� ��40 �2@� 0��� � ����3�/� �����K� ��� H-�����M� �� � �0K� �� �� ��D0 �2@� 0��� � ����3�/� �����K� ��� H-����H0 �2@� 0��3�/� ��� H-�����M� �� �p0 �2@� 0��3�/� �m����K� ��� H-�����M� �� �H0 �2@� 0��3�/��K� ����-� ����M� �0�(��  ��0�T �� �� ��?�2@�0��0�  �� ���3�2@�  ��0� ���3�2@�  ��0� ��0�$�  �� �< �0@�$0��0�  ��( �� 0�2@� 0��#8��  S�  $0�2@�  ��< �0@� R�   0�2@�  ��0�0 �� �S<�S9D�40��0�!��@ ��0�!��D �� � 0 ��?K�H0��0�&��L �� �S<�S9D�P0�� 0�� �� Ћ� ���/��-� ����M� �� �4 �0A�  ��  �� 4 �0A� ��  ��$4 �0A�  ��  ��(4 �0A�  ��  ��,4 �0A�  ��  ��0��0� 4 �0A� �  ��4 �0A� 0��0�0�0�  S�   0��Z  �04 �0A�   � A�  ��  ��44 �0A�  � A�  ��  ��84 �0A�  � A�  ��  ��<4 �0A�  � A�  ��  ��@4 �0A� �  ��4 �0A� 0��0�0�@0�  S����
4 �0A�@ ��  ��0�0� 5 �0A�  ��0�  ��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0�0�5 �0A�  ��0�  ��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0�� 0�� �� Ћ� ���/� H-����8�M�0 �4�8 �<0� K�(0K� ����  ��/O�h��� 0��  S�  
 0��K �2 �0A� 0��0�0�0�  S�  
 0��A �4 �0A� 0��0�0�0�  S�   0��7 �(0 �0A� ��  ��80 �0A� ��  ��0 �0A� ��  ��0��0�0�0��0�0�
=��0�0�;��0� 2 �0A� �  ��0��0�0�0��0�4 �0A� �  ��2 �0A� �  ��2 �0A� �  ��2 �0A� �  ��2 �0A� �  ��02 �0A�( �  ��42 �0A�$ �  ��82 �0A�  �  ��<2 �0A� �  ��p4 �0A� �  ��t4 �0A� �  ��x4 �0A� �  ��|4 �0A� �  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A� ��  �� 4 �0A�< �  ��$4 �0A�  ��  ��(4 �0A�  ��  ��,4 �0A�  ��  ��0��0� 4 �0A� �  ��00 �0A�4 �  ��40 �0A�< �  �� 0 �0A�0 �  ��$0 �0A�< �  ��0 �0A� 0��0�0�0�  S����
0 �0A� ��  ��2 �0A�  ��  ��2 �0A�  ��  ��2 �0A�  ��  ��2 �0A�  ��  ��02 �0A�  ��  ��42 �0A�  ��  ��82 �0A�  ��  ��<2 �0A�  ��  ��4 �0A� 0��0�0�@0�  S����
4 �0A�@ ��  ��p4 �0A�  ��  ��t4 �0A�  ��  ��x4 �0A�  ��  ��|4 �0A�  ��  ��80�  �� 5 �0A� 0�� R�9  80�0��  ��5 �0A� 0�� R�1  80�0��  ��5 �0A� 0�� R�)  80�0��  ��5 �0A� 0�� R�!  80�0��  ��5 �0A� 0�� R�  80�0��  ��5 �0A� 0�� R�  80�0��  ��5 �0A� 0�� R�	  80�0��  ��5 �0A� 0�� R�   0��   � 0�� ���K� ��� H-����8�M�8 � 0�2@�0�9��0�  K�00K� ����  ��/O���� 0��  S�  
 0���  �4 �0A� 0��0�0�0�  S�   0���  �0 �0A�  ��  ��p4 �0A�  �  ��t4 �0A� �  ��x4 �0A� �  ��|4 �0A� �  ��4 �0A�8 �  ��  ��4 �0A�8 � ��  ��  ��4 �0A�8 � ��  ��  ��4 �0A�8 � ��  ��  ��4 �0A�8 � ��  ��  ��4 �0A�8 � ��  ��  ��4 �0A�8 � ��  ��  ��4 �0A�8 � ��  ��  ��4 �0A� ��  �� 4 �0A� �  ��$4 �0A�  ��  ��(4 �0A�  ��  ��,4 �0A�  ��  ��0��0� 4 �0A� �  ��@0 �0A� �  ��D0 �0A� �  ��0 �0A� 0��0�  S����
0 �0A� ��  ��4 �0A� 0��0�0�@0�  S����
4 �0A�@ ��  ��p4 �0A�  ��  ��t4 �0A�  ��  ��x4 �0A�  ��  ��|4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  �� 5 �0A�  ��80�  ��80� ��5 �0A� 0�� 0��80� ��5 �0A� 0�� 0��80� ��5 �0A� 0�� 0��80� ��5 �0A� 0�� 0��80� ��5 �0A� 0�� 0��80� ��5 �0A� 0�� 0��80� ��5 �0A� 0�� 0�� 0�� ���K� ����-� ����M� �� �0�  S�   0��Z  �H0 �0A� ��  ��4 �0A� ��  ��0 �0A� 0��0�0�0��0�0 �0A� �  ��0��0� 4 �0A� �  ��4 �0A� ��  �� 4 �0A� �  ��$4 �0A�  ��  ��@0 �0A� �  ��D0 �0A� �  ��4 �0A� 0��@0�  S����
4 �0A�@ ��  ��0�0� 5 �0A�  ��0�  ��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0 �0A� ��  �� 0�� �� Ћ� ���/� H-����0�M�  �$�( �,0�(0� K� ��$� ����� 0�3>��,0�� 0����� 0� ��0K�,� ������ ��C�� ��0��<�/� 0��0�0� ���K� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ������������������ �À�����@�à�� ��xV4  ��� �= ���  � ��� �� �)�C  ��ӟ����  ��� � @��P��`��Р� O� P�#  
��\ �\0� �� �� �� P����:x � �Fఠ�� ��� ��  ���0�� 0��  ��	 �����p� W�  
 W�   
  �!������	��  � ��	�� �� �� R����:� ����0�@�� ����  ��  �� �� P���� ��VO���� ������4]  � 4{ 4{ �  �  �����
�� ��
�� ��������  ����� � � � � � � � �|�� ��� �O����Р��i�����H�M����!� ��H ��4P���� �� �� � � � � � � � � � � � � ��M�  ���� ���  O����  ��Ѝ�H�M����"� ��H ��4P���� �� ��t � � � � � � � � � � � � �<�� ��� �O����Р��i�����H�M����d"� ��H ��4P���� �� ��S � � � � � � � � � � � � ��� ��� �O����Р��i�����H�M�����"� ��H ��4P���� �� ��2 � � � � � � � � � � � � ���� ��� �O����Р��i�����H�M����$#� ��H ��4P���� �� �� � � � � � � � � � � � � �\�� ��� �O����Р��i�����H�M����#� ��H ��4P���� �� ��� � � � � � � � � � � � � ��� ��� �O����Р��i�����H�M�����#� ��H ��4P���� �� ��� �  �B � � � � � � � � � �  ��� �  �!(��0 R�0 �0���ӟ� @-� ����� ����� ����� ���#�� Q�?  
��� ���� ����� ��� ����� ����� �� ����� ���� �� ��� ��>  ��� ��� �  �� Q�  
�� ��!��� Q�  �  �] �  �[ �v �U  �  �  ��i �    5  �@��C/����9������  �(�� @� �� �� ������ ��  �� ��[��  ����� �� ���� ��!��� Q�  �2��$���  Q�   �  �1 �  �/ �J �\  �b ��� ��> � R�0� R�0� R�0�( R�0����0����E��|�� ��x��x�� ��t��t��t"����p��p"����<��h������ ��\����5��(����,��H�� �������� Q�  
 Q�  
 Q�  
 Q����
���"��������  ���� ������� ���� ���������� ��*�� Q��� @� 0��0�3 0�����:  � ����� �����������x��!�����������������, ����x!��x ��x �� P�����O��o���� � � � � � � ��  �                                         � � � ������ � ��  Q��/���� � ��P��_�� ����� �� ������ ��� � � � � � � � ��� ���0��\@��P��P��P�����#�� �� ��
����  ��	��  t��  3` h d � �    �C  �KKKK   """"  @"""   fff P�  www P�    �  OOOOH�  \ UL�   ���   ���  �� � � � � � �@�� ����
�� @-� R���� ��� @-��������$����������D�������������������������������������� �������������������x����]��0��l��4��h��8��d��<��d ����������*������H����',������<����?.������0��������$���� �����D��������������������������������������� �����������������������]��0����4��|��8��x��<��d ���������*�����\����',�����P����?.�����D��������8���� ��� @-���� �� �� ��$����D������������������������������������������� ���������������������������0��|����4����8����<��d ��P�������*��L�������',��H�������?.��D�����������?.��>���B����?.��:���
����?.��6������������ ����*��.�������������*��(������ �� �� ��$�����D��������������l��������������������L�� ������|�������������0������0��$��T��4��P��8��L��<��d ����������*����������',����������?.��������������?.������B����?.������
����?.�������������������*��������������*������@ �� ��  ��  ���� �� ��` �� ��  ��  ���� �� �� ���  w     `T��q
q�0� %  #�@� @���I436e8P  �       aU��   �    &0 3�@OeFx@F<
 Rq�� Q������������
��@�� ����
�� @-��� �� #����Q+���2����������"��������"���� ���"�����"���2������ ���"�����"���2����������"������B,����+��!0��������E,������,����!+��!0��������,������)����|��|"����x��x"����t��t"����p��p"����l��l"����h��h"����d��d"����`"����\2�� Q�  <��P"����L��<"������@"����<��<"����8��8"������0"������("����$��$"�����!������!������!�����"����� ��X!����Q+���1��������!����A+���1��{�����@!����<!���1��u�����4!����0!��1��o����� ��!��� Q�8  �1��$���  Q�3  ����� ������ ������ ����a����� ������ ����Z���X��H�� ����@�� ����8�� ����O����� ������ ����H��� ����  ���� �� ��  ����� ����� ����� ����� ���� ���   B      �  �  �  �  tT!�  *    p  �  (#   �    E   E  8  A  }� A  d�  d��    f�  @��  (�  $�  �� �       !!!    `
�  �  a�0�3%    ���/� ��"���N-� ��� ����M� ���  �� p�� �� ��  �� `�� �� ��  �� P��$ �� ��  �� @��, �� ��  �� ���4 �� ��  ��< ��D ��  ��  �� 0��L ����L �� ��#��`��&B�L ��  ���� ������ ���� ��(���� ��0���� ��8���� ��@����  ��H��Ѝ�����D ��1��s����/�@-�� � �(0�� 0��0C� S�  �Ho �l �  �l �Do �  ��������@-�0��8�� S�   ����J< �  �����  N��V��  ����tr ��@-��M� ��	 �� ��[� �� �� �� ��a �0��w S�0   ����� ��Z � ��"��� ��V � ��+��� ��R � ����� ��N � ��!��� ��J � ��*��� ��F � ��H��� ��B ������>C �����;C �����8C �����5C �����2C �����/C �����X  � S�p��`��P��@��  � ��3��� ��# � ��5��� �� � ��>��� �� � ��G��� �� ���0��C �����C ��� ��C ������6  � ���� �� � ���� �� � ��(�� ��� � ���� ��� ��� �� ��� � �� �� ��� ��� �� ��� � ��&�� ��� ���d���B ���\���B ���T���B ���\���B ���@���B ���8���B ���0���B �4����@���B �(���B �$�� �� ��� ������B �1��P3�� S�  ���B � ��$���������0��� ��@�� ��"��@�������������������(B� ���  �� �����������(���� �������� �����  ��B � 0�� S� �  
S� �  
 S� �  
 S�| �  
 S�  p ��B �  ��Ѝ�����������������
����*��:��G��W���n��  ��""""  "   W���  @��������������������/�E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� �����E5��$ �� ��$ ��$ �� ��$ �����E5��$ �� ��$ ��$ �� ��$ �����E5��$ �� ��$ ��$ �� ��$ �����E5��$ �� ��$ ��$ �� ��$ �����@-����������@�����@-����������@�����@-�����������@������@-����������@�����@-�������������@������@-�����������@������@-�y������v���@�����@-����z���p���@��o���@-�EE���0��0���0���0��0���0��e����0��0���0��a����0���0��0���0��\����0��0���0��X����0��0��0���0��@��k���E5��� �� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��S���@-�Y���`���6���@��m���@-�k���Z���0���@��O���@-�EE���0��<���0���0��0���0��%����0��0���0��!����0���0��0���0������0��0���0������0��<��<���0��@��K���@-�Q���X������@��e���@-�c���R������@��G���@-�EE�� 0��<�� 0��$0��0��$0������$0��0��$0������$0��$0��0��$0������$0��0��$0������ 0��<��<�� 0��@��C���E5��� �� ��� ��� �� ��� ��� �� ��� ��� ��� �� ��� ��� �� �� ��� ������E5��� ��� ��� ��� �� ��� ��� �� ��� ��� ��*��*��� ��� ��,��,��� ������E5��( ��� ��( ��$ �� ��$ ��$ �� ��$ ��  ��*��*��  ��  ��,��,��  ������A-� @��P��p��1���`��T6�� �  
���   ����`V�������@��1���@D�U4�� �  
���   �����  T����'���@��@D�W4�� �  
����   �����  T��������A������D-� @��P��p��	���`��T6�� �  
����   �����`V��������`��	���`F�U6�� �  
����   �����  V��������P������T5�� �  
����   �����PU��������`������E5��� �� ��� ��� �� ��� ��� �� ��� ��V���EE��`F��0��0���0���0��0���0��M����0��0���0���0��0���0��F���Ġ���0���
�0���0���0��V��0���0��<����0��uP��0���0���0��0���0��4���  V���������0��0��0���0����� P�������A-� @��P��p������`��T6�� �  
����   ����`V��������@������@D�U4�� �  
����   ����  T��������@��@D�W4�� �  
|���   �t���  T���������A�������A-� @��P��p������`��T6�� �  
w���   �o���`V����l���@������@D�U4�� �  
k���   �c���  T��������@��@D�W4�� �  
`���   �X���  T���������A������s@-� @P�`��  
 T� @�!P�  
 T� @�*P�  
 T� @�,P�	  
 T�@�HP�  
 T�@�DP�  
����P���� ��� ��2���0�� ����$��� ��D��t �� �����|����@-� PP�p��`��  
 U�"@�  
 U�+@�
  
 U�-@�  
 U�H@�  
 U�D@�  
����@���� ��� ��?p���� ����� ��? �� �� ������ �����������  P� ��  
 P�5�
  
 P�>�  
 P�G�  
 P�P�  
����3��� ������4��`,��*��`,��d,�� ��d,���/�4��`,��*��`,��d,��  ��d,���/�p `��/� P�0@-�  1��? �� ��).�� ��X �� ��  � Q� Q1�).� �8 � �0P����� @�� ��0��� �� P��P��@��P��RZ��P��0@������  �C L P�@-�  1���" � ��N/�� ��X �� ��  � Q� Q1�N/� �8 � �0@����� ��� ��$0�� @��'J��@��@��@�� @��@��@����� �  �C L ��� �� �� 0�����  ��� �� ��0������ �� ��p `� ���/�@-�? ��)�� ��0����0�����  �C  @-�0����p�����  @-�)����0����4�����  �C  @-���0��)����D�����  �C  @-�0����H�����    ��p@-� P��@��0��@����  T� ����� ��� ��`��0�� ��<��@ ��c �`��p�������� 0��  �� ����~c ������ 0��  �� �����c �����6�� ��@-� �� ��@�� �� �� �� �� �� ��  �� �� �� ��0��0��0��  ��6��  ��@�����@��@�� �� �� ����� �� ��0 �� ���6��(0�� ����
 0���&��������0��S����0������0��0��Q����  �����  �C� ���/� ���/�@-�@��p ��T��A������  ��H������D��t ��������8������  ��0������  ��(������0��8�� ����
��� ��� ���@�@-� ������0����C3C� P� ����  @-� @�� ��������(0��  �S�����0�� �� S�+B�#B�������   p@-�H`��@�� P�� �� ����@������@ T�k��  P�� ������ @P����0�� V����p���  �C  �C@-�  ��> �0�� �� $��~T �  P����
@��jT ����  0��$��  ���/����$0��P����@-� 0��@�� �������� ��������0��P�� 0�� ���/����$0��P�� ��@-� 0��@�� �������� ��������0��P�� �� 0�� ���/����0��P�� �� 0�� ��P��  ��/����0��P�� �� 0�� ���/����(0��P�� ����@-� 0��@�� �������� ��������0��P�� �� 0�� ���/����$0��P����@-� 0��@�� �������� ��������0��P�� 0�� ���/����(0��P�� ����@-� 0��@�� �������� �������� 0��P�� ��  �� 1��#8��8��0�� 1���/����0��P�� �� 0�� ���/����0��P�� �� 0�� ���/���� ��0��0�� �� ��0���/���� 
@  �����0��  ���������/���� 	@  ��0�� �� �� �� ��  ��  �� ���/� 	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/���� 
@  �����0��  ���������/���� 	@  ��0�� �� �� �� ��  ��  �� ���/� 	@ ��� ��0��0�� �� ��0���/����$
@  �����0��  ���������/����$	@  ��0�� �� �� �� ��  ��  �� ���/�$	@ ��� ��0��0�� �� ��0���/����(
@  �����0��  ���������/����(	@  ��0�� �� �� �� ��  ��  �� ���/�(	@ ��� ��0��0�� �� ��0���/����,
@  �����0��  ���������/����,	@  ��0�� �� �� �� ��  ��  �� ���/�,	@ ��� ��0��0�� �� ��0���/����0
@  �����0��  ���������/����0	@  ��0�� �� �� �� ��  ��  �� ���/�0	@ ��� ��0��0�� �� ��0���/����4
@  �����0��  ���������/����4	@  ��0�� �� �� �� ��  ��  �� ���/�4	@ ��� ��0��0�� �� ��0���/����8
@  �����0��  ���������/����8	@  ��0�� �� �� �� ��  ��  �� ���/�8	@ ��� ��0��0�� �� ��0���/����<
@  �����0��  ���������/����<	@  ��0�� �� �� �� ��  ��  �� ���/�<	@ ��� ��0��0��  �� :���/����0���� 0�� )�� �� )���/����0�� ��0��  �� 9�� 0��  �� 	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  �� :���/����0���� 0�� )�� �� )���/����0�� ��0��  �� 9�� 0��  �� 	���/���� ��0��0��  ��@?���/����0���� 0�� /�� �� /���/����0�� ��0��  �� ?�� 0��  �� ���/���� ��0��0��  ��D?���/����0���� 0��/�� ��/���/����0�� ��0��  ��?�� 0��  �����/���� ��0��0��  ��H?���/����0���� 0��/�� ��/���/����0�� ��0��  ��?�� 0��  �����/���� ��0��0��  ��L?���/����0���� 0��/�� ��/���/����0�� ��0��  ��?�� 0��  �����/���� ��0��  �����������/���� @ 0�� 0�� +�� �� �� +���/���� �� @� �� ��0��  ���� ��  �� ���/����@ 0�� @� ��0�� 0��+��  ��  �����/����0��  ��0�� ���/����@ 0�� 0�����/����0��  ��0�� ���/����@ 0�� 0�����/���� ��0��  �����������/����@ 0�� 0��+�� �� ��+���/����0@� S�	  �(0�� @� 0��>��0�� !�� ���� ���/� ��: ������ @� P�o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ������������������ �À�����@�à�� ��xV4  ��� �= ���  � ��� �� �)�C  ��ӟ����  ��� � @��P��`��Р� O� P�#  
��\ �\0� �� �� �� P����:x � �Fఠ�� ��� ��  ���0�� 0��  ��	 �����p� W�  
 W�   
  �!������	��  � ��	�� �� �� R����:� ����0�@�� ����  ��  �� �� P���� ��VO���� ������4]  � 4{ 4{ �  �  �����
�� ��
�� ��������  ����� � � � � � � � �|�� ��� �O����Р��i�����H�M����!� ��H ��4P���� �� �� � � � � � � � � � � � � ��M�  ���� ���  O����  ��Ѝ�H�M����"� ��H ��4P���� �� ��t � � � � � � � � � � � � �<�� ��� �O����Р��i�����H�M����d"� ��H ��4P���� �� ��S � � � � � � � � � � � � ��� ��� �O����Р��i�����H�M�����"� ��H ��4P���� �� ��2 � � � � � � � � � � � � ���� ��� �O����Р��i�����H�M����$#� ��H ��4P���� �� �� � � � � � � � � � � � � �\�� ��� �O����Р��i�����H�M����#� ��H ��4P���� �� ��� � � � � � � � � � � � � ��� ��� �O����Р��i�����H�M�����#� ��H ��4P���� �� ��� �  �B � � � � � � � � � �  ��� �  �!(��0 R�0 �0���ӟ� @-� ����� ����� ����� ���#�� Q�?  
��� ���� ����� ��� ����� ����� �� ����� ���� �� ��� ��>  ��� ��� �  �� Q�  
�� ��!��� Q�  �  �] �  �[ �v �U  �  �  ��i �    5  �@��C/����9������  �(�� @� �� �� ������ ��  �� ��[��  ����� �� ���� ��!��� Q�  �2��$���  Q�   �  �1 �  �/ �J �\  �b ��� ��> � R�0� R�0� R�0�( R�0����0����E��|�� ��x��x�� ��t��t��t"����p��p"����<��h������ ��\����5��(����,��H�� �������� Q�  
 Q�  
 Q�  
 Q����
���"��������  ���� ������� ���� ���������� ��*�� Q��� @� 0��0�3 0�����:  � ����� �����������x��!�����������������, ����x!��x ��x �� P�����O��o���� � � � � � � ��  �                                         � � � ������ � ��  Q��/���� � ��P��_�� ����� �� ������ ��� � � � � � � � ��� ���0��\@��P��P��P�����#�� �� ��
����  ��	��  t��  3` h d � �    �C  �KKKK   """"  @"""   fff P�  www P�    �  OOOOH�  \ UL�   ���   ���  �� � � � � � �@�� ����
�� @-� R���� ��� @-��������$����������D�������������������������������������� �������������������x����]��0��l��4��h��8��d��<��d ����������*������H����',������<����?.������0��������$���� �����D��������������������������������������� �����������������������]��0����4��|��8��x��<��d ���������*�����\����',�����P����?.�����D��������8���� ��� @-���� �� �� ��$����D������������������������������������������� ���������������������������0��|����4����8����<��d ��P�������*��L�������',��H�������?.��D�����������?.��>���B����?.��:���
����?.��6������������ ����*��.�������������*��(������ �� �� ��$�����D��������������l��������������������L�� ������|�������������0������0��$��T��4��P��8��L��<��d ����������*����������',����������?.��������������?.������B����?.������
����?.�������������������*��������������*������@ �� ��  ��  ���� �� ��` �� ��  ��  ���� �� �� ���  w     `T��q
q�0� %  #�@� @���I436e8P  �       aU��   �    &0 3�@OeFx@F<
 Rq�� Q������������
��@�� ����
�� @-��� �� #����Q+���2����������"��������"���� ���"�����"���2������ ���"�����"���2����������"������B,����+��!0��������E,������,����!+��!0��������,������)����|��|"����x��x"����t��t"����p��p"����l��l"����h��h"����d��d"����`"����\2�� Q�  <��P"����L��<"������@"����<��<"����8��8"������0"������("����$��$"�����!������!������!�����"����� ��X!����Q+���1��������!����A+���1��{�����@!����<!���1��u�����4!����0!��1��o����� ��!��� Q�8  �1��$���  Q�3  ����� ������ ������ ����a����� ������ ����Z���X��H�� ����@�� ����8�� ����O����� ������ ����H��� ����  ���� �� ��  ����� ����� ����� ����� ���� ���   B      �  �  �  �  tT!�  *    p  �  (#   �    E   E  8  A  }� A  d�  d��    f�  @��  (�  $�  �� �       !!!    `
�  �  a�0�3%    ���/� ��"���N-� ��� ����M� ���  �� p�� �� ��  �� `�� �� ��  �� P��$ �� ��  �� @��, �� ��  �� ���4 �� ��  ��< ��D ��  ��  �� 0��L ����L �� ��#��`��&B�L ��  ���� ������ ���� ��(���� ��0���� ��8���� ��@����  ��H��Ѝ�����D ��1��s����/�@-�� � �(0�� 0��0C� S�  �Ho �l �  �l �Do �  ��������@-�0��8�� S�   ����J< �  �����  N��V��  ����tr ��@-��M� ��	 �� ��[� �� �� �� ��a �0��w S�0   ����� ��Z � ��"��� ��V � ��+��� ��R � ����� ��N � ��!��� ��J � ��*��� ��F � ��H��� ��B ������>C �����;C �����8C �����5C �����2C �����/C �����X  � S�p��`��P��@��  � ��3��� ��# � ��5��� �� � ��>��� �� � ��G��� �� ���0��C �����C ��� ��C ������6  � ���� �� � ���� �� � ��(�� ��� � ���� ��� ��� �� ��� � �� �� ��� ��� �� ��� � ��&�� ��� ���d���B ���\���B ���T���B ���\���B ���@���B ���8���B ���0���B �4����@���B �(���B �$�� �� ��� ������B �1��P3�� S�  ���B � ��$���������0��� ��@�� ��"��@�������������������(B� ���  �� �����������(���� �������� �����  ��B � 0�� S� �  
S� �  
 S� �  
 S�| �  
 S�  p ��B �  ��Ѝ�����������������
����*��:��G��W���n��  ��""""  "   W���  @��������������������/�E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� ������E5��� �� ��� ��� �� ��� �����E5��$ �� ��$ ��$ �� ��$ �����E5��$ �� ��$ ��$ �� ��$ �����E5��$ �� ��$ ��$ �� ��$ �����E5��$ �� ��$ ��$ �� ��$ �����@-����������@�����@-����������@�����@-�����������@������@-����������@�����@-�������������@������@-�����������@������@-�y������v���@�����@-����z���p���@��o���@-�EE���0��0���0���0��0���0��e����0��0���0��a����0���0��0���0��\����0��0���0��X����0��0��0���0��@��k���E5��� �� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��� �� ��� ��S���@-�Y���`���6���@��m���@-�k���Z���0���@��O���@-�EE���0��<���0���0��0���0��%����0��0���0��!����0���0��0���0������0��0���0������0��<��<���0��@��K���@-�Q���X������@��e���@-�c���R������@��G���@-�EE�� 0��<�� 0��$0��0��$0������$0��0��$0������$0��$0��0��$0������$0��0��$0������ 0��<��<�� 0��@��C���E5��� �� ��� ��� �� ��� ��� �� ��� ��� ��� �� ��� ��� �� �� ��� ������E5��� ��� ��� ��� �� ��� ��� �� ��� ��� ��*��*��� ��� ��,��,��� ������E5��( ��� ��( ��$ �� ��$ ��$ �� ��$ ��  ��*��*��  ��  ��,��,��  ������A-� @��P��p��1���`��T6�� �  
���   ����`V�������@��1���@D�U4�� �  
���   �����  T����'���@��@D�W4�� �  
����   �����  T��������A������D-� @��P��p��	���`��T6�� �  
����   �����`V��������`��	���`F�U6�� �  
����   �����  V��������P������T5�� �  
����   �����PU��������`������E5��� �� ��� ��� �� ��� ��� �� ��� ��V���EE��`F��0��0���0���0��0���0��M����0��0���0���0��0���0��F���Ġ���0���
�0���0���0��V��0���0��<����0��uP��0���0���0��0���0��4���  V���������0��0��0���0����� P�������A-� @��P��p������`��T6�� �  
����   ����`V��������@������@D�U4�� �  
����   ����  T��������@��@D�W4�� �  
|���   �t���  T���������A�������A-� @��P��p������`��T6�� �  
w���   �o���`V����l���@������@D�U4�� �  
k���   �c���  T��������@��@D�W4�� �  
`���   �X���  T���������A������s@-� @P�`��  
 T� @�!P�  
 T� @�*P�  
 T� @�,P�	  
 T�@�HP�  
 T�@�DP�  
����P���� ��� ��2���0�� ����$��� ��D��t �� �����|����@-� PP�p��`��  
 U�"@�  
 U�+@�
  
 U�-@�  
 U�H@�  
 U�D@�  
����@���� ��� ��?p���� ����� ��? �� �� ������ �����������  P� ��  
 P�5�
  
 P�>�  
 P�G�  
 P�P�  
����3��� ������4��`,��*��`,��d,�� ��d,���/�4��`,��*��`,��d,��  ��d,���/�p `��/� P�0@-�  1��? �� ��).�� ��X �� ��  � Q� Q1�).� �8 � �0P����� @�� ��0��� �� P��P��@��P��RZ��P��0@������  �C L P�@-�  1���" � ��N/�� ��X �� ��  � Q� Q1�N/� �8 � �0@����� ��� ��$0�� @��'J��@��@��@�� @��@��@����� �  �C L ��� �� �� 0�����  ��� �� ��0������ �� ��p `� ���/�@-�? ��)�� ��0����0�����  �C  @-�0����p�����  @-�)����0����4�����  �C  @-���0��)����D�����  �C  @-�0����H�����    ��p@-� P��@��0��@����  T� ����� ��� ��`��0�� ��<��@ ��c �`��p�������� 0��  �� ����~c ������ 0��  �� �����c �����6�� ��@-� �� ��@�� �� �� �� �� �� ��  �� �� �� ��0��0��0��  ��6��  ��@�����@��@�� �� �� ����� �� ��0 �� ���6��(0�� ����
 0���&��������0��S����0������0��0��Q����  �����  �C� ���/� ���/�@-�@��p ��T��A������  ��H������D��t ��������8������  ��0������  ��(������0��8�� ����
��� ��� ���@�@-� ������0����C3C� P� ����  @-� @�� ��������(0��  �S�����0�� �� S�+B�#B�������   p@-�H`��@�� P�� �� ����@������@ T�k��  P�� ������ @P����0�� V����p���  �C  �C@-�  ��> �0�� �� $��~T �  P����
@��jT ����  0��$��  ���/����$0��P����@-� 0��@�� �������� ��������0��P�� 0�� ���/����$0��P�� ��@-� 0��@�� �������� ��������0��P�� �� 0�� ���/����0��P�� �� 0�� ��P��  ��/����0��P�� �� 0�� ���/����(0��P�� ����@-� 0��@�� �������� ��������0��P�� �� 0�� ���/����$0��P����@-� 0��@�� �������� ��������0��P�� 0�� ���/����(0��P�� ����@-� 0��@�� �������� �������� 0��P�� ��  �� 1��#8��8��0�� 1���/����0��P�� �� 0�� ���/����0��P�� �� 0�� ���/���� ��0��0�� �� ��0���/���� 
@  �����0��  ���������/���� 	@  ��0�� �� �� �� ��  ��  �� ���/� 	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/����
@  �����0��  ���������/����	@  ��0�� �� �� �� ��  ��  �� ���/�	@ ��� ��0��0�� �� ��0���/���� 
@  �����0��  ���������/���� 	@  ��0�� �� �� �� ��  ��  �� ���/� 	@ ��� ��0��0�� �� ��0���/����$
@  �����0��  ���������/����$	@  ��0�� �� �� �� ��  ��  �� ���/�$	@ ��� ��0��0�� �� ��0���/����(
@  �����0��  ���������/����(	@  ��0�� �� �� �� ��  ��  �� ���/�(	@ ��� ��0��0�� �� ��0���/����,
@  �����0��  ���������/����,	@  ��0�� �� �� �� ��  ��  �� ���/�,	@ ��� ��0��0�� �� ��0���/����0
@  �����0��  ���������/����0	@  ��0�� �� �� �� ��  ��  �� ���/�0	@ ��� ��0��0�� �� ��0���/����4
@  �����0��  ���������/����4	@  ��0�� �� �� �� ��  ��  �� ���/�4	@ ��� ��0��0�� �� ��0���/����8
@  �����0��  ���������/����8	@  ��0�� �� �� �� ��  ��  �� ���/�8	@ ��� ��0��0�� �� ��0���/����<
@  �����0��  ���������/����<	@  ��0�� �� �� �� ��  ��  �� ���/�<	@ ��� ��0��0��  �� :���/����0���� 0�� )�� �� )���/����0�� ��0��  �� 9�� 0��  �� 	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  ��:���/����0���� 0��)�� ��)���/����0�� ��0��  ��9�� 0��  ��	���/���� ��0��0��  �� :���/����0���� 0�� )�� �� )���/����0�� ��0��  �� 9�� 0��  �� 	���/���� ��0��0��  ��@?���/����0���� 0�� /�� �� /���/����0�� ��0��  �� ?�� 0��  �� ���/���� ��0��0��  ��D?���/����0���� 0��/�� ��/���/����0�� ��0��  ��?�� 0��  �����/���� ��0��0��  ��H?���/����0���� 0��/�� ��/���/����0�� ��0��  ��?�� 0��  �����/���� ��0��0��  ��L?���/����0���� 0��/�� ��/���/����0�� ��0��  ��?�� 0��  �����/���� ��0��  �����������/���� @ 0�� 0�� +�� �� �� +���/���� �� @� �� ��0��  ���� ��  �� ���/����@ 0�� @� ��0�� 0��+��  ��  �����/����0��  ��0�� ���/����@ 0�� 0�����/����0��  ��0�� ���/����@ 0�� 0�����/���� ��0��  �����������/����@ 0�� 0��+�� �� ��+���/����0@� S�	  �(0�� @� 0��>��0�� !�� ���� ���/� ��: ������ @� P�  �$ ��$0��  ��0�� !�� ���� ���/� ��r: ����@ ��0������0��P�� 0�� !�� ���� ���/�����D-�p���0�� P� @��P��`�� ���  ڼ ��X: � W�  ڰ ��T: � T�  ʤ0��!��������������R��P������ T�  �h ��A��p0��������  �� ����D��a��`������@D� T������A��<0�� ��� ��b�� ��t��  ����D��@��@�����������%�� @  @ @ �D-�p���0�� P�`�� @��$��P��  ��  �� ��: � W�  ڴ ��: � T�  ʨ0��$�������� ����������\��P����� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��@   @ @ @ �D-�p���0�� P�`�� @��$��P��  ��  �� ���9 � W�  ڴ ���9 � T�  ʨ0��$�������� ����������\��P��U��� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��@ @ @ @ @ �D-�p��0�� P�`�� @��$��P��  ��  ڠ ��9 � W�  ڔ ��9 � T����Ȉ0��$��������| ����������\��P����� T�L0��
  
  ��A��P0�������� ����D��a��`������  ��,0�������c��p��p�����������%��@ ` @ @ @ �D-�p��0�� P�`�� @��$��P��  ��  ڠ ��Z9 � W�  ڔ ��V9 � T����Ȉ0��$��������| ����������\��P������ T�L0��
  
  ��A��P0�������� ����D��a��`������  ��,0�������c��p��p�����������%��@ � @  @ $@ �D-�p��0�� P�`�� @��$��P��  ��  �x �� 9 � W�  �l ��9 � T�����`0��$����������P �����A�����\��P�����$ ��40��������  �� ����D��a��`�����������%��@ � @ (@ �D-�p��0�� P�`�� @��$��P��  ��  �x ���8 � W�  �l ���8 � T�����`0��$����������P �����A�����\��P��o���$ ��40��������  �� ����D��a��`�����������%��@ � @ 0@ �D-�p��0�� P�`�� @��$��P��  ��  ڠ ���8 � W�  ڔ ��8 � T����Ȉ0��$��������| ����������\��P��A��� T�L0��
  
  ��A��P0�������� ����D��a��`������  ��,0�������c��p��p�����������%��@ � @ 8@ <@ �D-�p���0�� P�`�� @��$��P��  ��  �� ��8 � W�  ڴ ��8 � T�  ʨ0��$�������� ����������\��P����� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%�� @  @ @@ D@ �D-�p���0�� P�`�� @��$��P��  ��  �� ��F8 � W�  ڴ ��B8 � T�  ʨ0��$�������� ����������\��P������ T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��$@  @ H@ L@ �D-�p���0�� P�`�� @��$��P��  ��  �� ��8 � W�  ڴ �� 8 � T�  ʨ0��$�������� ����������\��P����� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��(@ @@ P@ T@ �D-�p���0�� P�`�� @��$��P��  ��  �� ���7 � W�  ڴ ��7 � T�  ʨ0��$�������� ����������\��P��A��� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��,@ `@ X@ \@ �D-�p���0�� P�`�� @��$��P��  ��  �� ��7 � W�  ڴ ��|7 � T�  ʨ0��$�������� ����������\��P������ T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��0@ �@ `@ d@ �D-�p���0�� P�`�� @��$��P��  ��  �� ��>7 � W�  ڴ ��:7 � T�  ʨ0��$�������� ����������\��P����� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��4@ �@ h@ l@ �D-�p���0�� P�`�� @��$��P��  ��  �� ���6 � W�  ڴ ���6 � T�  ʨ0��$�������� ����������\��P��{��� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��8@ �@ p@ t@ �D-�p���0�� P�`�� @��$��P��  ��  �� ��6 � W�  ڴ ��6 � T�  ʨ0��$�������� ����������\��P��9��� T�  �h ��A��t0��������  �� ����D��a��`������@D� T������A��@0�� ��� ��b�� ��t��  ����D��@��@�����������%��<@ �@ x@ |@ �@-�p���0�� P�`�� @��$��P��  ��  ڴ ��x6 � W�  ڨ ��t6 � T�  �4��!�� Ǔ���  �������R�� W������ T�
  �`0��A��� �� �� 0�� ����D��b�� h������@D� T������A�����0��c��0��t�� 0��(��D��@��H�����������%���@-�p��0�� P�`�� @��$��P��  ��  ڔ ��=6 � W�  ڈ ��96 � T�����4��!��Ǔ���  �������R��W����� T�D0��	  
 0��A��� �� ������D��b��h������ 0��(��� ��c��p��x�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��
6 � W�  ڨ ��6 � T�  �4��!��Ǔ���@ �������R��W����� T�
  �`0��A��� �� �� 0������D��b��h������@D� T������A�����0��c��0��t�� 0��(��D��@��H�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ���5 � W�  ڨ ���5 � T�  �4��!��Ǔ���` �������R��W��O��� T�
  �`0��A��� �� �� 0������D��b��h������@D� T������A�����0��c��0��t�� 0��(��D��@��H�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��5 � W�  ڨ ��5 � T�  �4��!��Ǔ��� �������R��W����� T�
  �`0��A��� �� �� 0�� ����D��b�� h������@D� T������A�����0��c��0��t�� 0��$(��D��@��$H�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��Y5 � W�  ڨ ��U5 � T�  �4��!��Ǔ��� �������R��W������ T�
  �`0��A��� �� �� 0��(����D��b��(h������@D� T������A�����0��c��0��t�� 0��,(��D��@��,H�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��5 � W�  ڨ ��5 � T�  �4��!��Ǔ���� �������R��W����� T�
  �`0��A��� �� �� 0��0����D��b��0h������@D� T������A�����0��c��0��t�� 0��4(��D��@��4H�����������%���@-�p��0�� P�`�� @��$��P��  ��  �p ���4 � W�  �d ���4 � T�����4��!��Ǔ������ �����A��R��W��b��� 0��� �� �� 0��8����D��b��8h�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��4 � W�  ڨ ��4 � T�  �4��!�� Ǔ����������R�� W��9��� T�
  �`0��A��� �� �� 0��@����D��b��@h������@D� T������A�����0��c��0��t�� 0��D(��D��@��DH�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��~4 �? W�  ڨ ��z4 � T�  �4��!�� Γ����������R�� ^������ T�
  �`0��A��� �� �� 0������D��b��n������@D� T������A�����0��c��0��t�� 0��.��D��@��N�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��C4 �? W�  ڨ ��?4 � T�  �4��!��Γ�����������R��^������ T�
  �`0��A��� �� �� 0������D��b��n������@D� T������A�����0��c��0��t�� 0��.��D��@��N�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ��4 �? W�  ڨ ��4 � T�  �4��!��Γ���1�������R��^����� T�
  �`0��A��� �� �� 0������D��b��n������@D� T������A�����0��c��0��t�� 0��.��D��@��N�����������%���@-�p���0�� P�`�� @��$��P��  ��  ڴ ���3 �? W�  ڨ ���3 � T�  �4��!��Γ�����������R��^��M��� T�
  �`0��A��� �� �� 0������D��b��n������@D� T������A�����0��c��0��t�� 0��.��D��@��N�����������%���@-�A��P���� �� `��9��`�� 0�屇 ���, ��(`��0��P�� p�� 0��;��$0�姇 �0��L ��t�� ��0��H ��<0��i��@p��D`�圇 �<0��l ��L��).��0��` ��\0��R:��d0��0��h0�吇 �\0�� �� ��N/��)>�� ��|0��':��0��	0��0�儇 �|0�� �����p��N?��`��0��0��0��z� �  U����*��0�0��0��@��� ��0��� ��&�� 0��� ��0�� ��� ��i� �0��� ����*��:��� ���0��6���0��0���0��]� �0��C��d��  ��0�� !���0��9��1��0��1��Q� ��0��  ���� �� @�� T�����������;��M��S��a��h���b��v��}�Á��0��  ���/�$ ��8@-�D ��3 �*  � @��&  �4�� P�� ��*� �$�� @�� ��&� ���  �� ��3 �  ��8�����@B ����/�  P�@-�80� 1�  
 P�	  (0��1��S��SH��0� ���ኣ �  ����_ � @   6n ������  ������0���� ��L��H%��D%���/� �  ` ��4���/��� ��P �� ���� �� ����<��@��H ��*�L ��, ��` ���-��h ��U-B�l �� ��0�� ���/�""" 03333 @D    U0��(��p@-� `�� ��x ��(��P�� Q�@��Q��\��  �A��Y��E��I��@��  �D0��D ��0�� S�  �80��Y��Y��0�I��@��  �  ��2 �0��P��@��p���?x}�����������@-��0�� @��@"��He��,��,��@"������奣 � p��P�� ����� �2 P�  ��0���l��`��`��He��  � U�@�����d0�� @��@"��Le��(��(��@"�����H�勣 � p��P�� ����� �P�  � 0���l��`��d��Le������ U�@��������� �@B X0���D-����He��k��� @��`���� � p��P�� ����� �
 P�  �0��D��HE������U�@��������� �@-�R �G �D � 0��?�?�S���  ����� P�����/� ���@-� @��B��A��A�� @����� ���@-� @����� @� T�   ����� \����  �����\ ����X0��Ƞ��  �� ��0@-� ���8 �� @�� P��@� ��, �� �������@����F�� ��ƌ� ��� @��0���  � ����0��  �� �� ���/���� ��  ��0�� ��  ��� �� ���/�@ ��������X0��X ���@-���  �� Q�  :�@��b�`��  �  ���@��  ��  b� `�� p�� ����� ��0�� �� ���������@ �@-� @������  d���� ���P�p@-� @�� �� @��	  :���P��d� �
�� `�� �`� ���  �  �����
�� �X� �<��V� � P��  ������@��0��  S�  *����@����� P����:p���< ����@B @-�  ������ ���������/��/��/��/��/��/��/��/��/��/� ����  �� ��80��0���/�@-��� ��1 �  �����\���	�� ��~1 �����	��<��� ��x �� ��P�၆ �(!��  ��< ��  �4�/�P��  P�   
����1��@��  T����8���A��� ���Ō�� ���Ɍ��P��,Ƞ�Ƞ�L���<0��q1 �� ��P��� ��  ��l1 �x�� ��� ��h1 �@P��  ��0�� 0����� ��0�� �� ��  �  ����0�� �� @�� S������ ��A1 � �� ��t ��� �p ��p@��x ��lP��  ���`�����4@��DP��H ��( ��b� �T��� �� ��������  �BH ��( �� ���5	��8��ð���[	�É	��D �ø	�Ëd��@ ��  ��0��ü0�� ��� @��P��  ��0��0��0��0��  �����A��A	E�o2 � ���X �@7 � �� @��( �ф � ��G �7 � �  �` ��( �  P�  
 �� ���� �H0��  ��D ��( � P�  
8 �� �㲗 ����, ���0 �  ��ٖ �]E �����D ������	���	��H ���	��4���	���N-� `�� ������������@��p��( � Z�  Z ���� P��p  ���w( �  P�  

�� �㲆 � p�� �����0 �	 ���� ��0��d��� ���h�������@ �  P�  
x���0 � ��WA �0��h�� ��`��� ������� �� ����  �� ����<1�� 0��  ���0������������ \������� �� ������ 1��  U� ���    �P�� 0��  S����
  S�  
�0�� ��̐��0��� �  ����0�� ��#1�� 0�嶄 � 0��  ��1�� 0��d ��  R�  
h0��  S�
  
|���b� 0�� �����p��� ��  �������� ���P0��  ��T �� 0��  �� ��}0 �2��� �������� ����� �������	���	���	��
�� ATD �� AT���	 AT BT-
�� ���  ����0��A� �� �� a�y� ��/���/���/��M� 0��  �  ��0��0��0��0��c S�����Ѝ��/� P�p@-� @��(  L����� 0��*���.�� ��!��0��
S����  ��L ����� 0��Q���1��P��P��#:��%Z����  ����� � S�ʠ��Ό�0�� �����: �� R������ 0��?����� P������ ���������� P������ ��p@�����
������@-����P����� ������@-����P����� P�p@-� @��  ���� �p��  �� �����@����� P����� ��p@����� ������
������0��  ��@ �� ��  ���/�L ���/�  ���/�p@-��M� @���� �� ��	� �0���,���<��8 ��40��� �� ������@P���/ �(��$ ��b� 0��� ���/ ������ ��0�� �� ����/ � ����� ��0�� �� ����/ �� ��Z �z ��C0�c0��V��v��  V� ���N��n���/ �@���T���@��P �� �0�H ����@ �1�� �4���0� ���/ �Ѝ�p������D
�É
�í
���
����V��·����a2��@-� ��=� �  ��@������<��@-� @�� ��/ � �����@������T��@-� @�� ��/ � �����@������O��@-� @�� ��/ � �����@������g��@-� @�� ��|/ � �����@������q��@-� @�� ��s/ � ��~���@������}��@-� @�� ��j/ � ��u���@��������@-� @�� ��a/ � ��l���@�������@-� ��E/ �P�� �a���  �����  ������� �� ��  ��M/ ���@-� @��� �� `����P������� ����  ������ ��������� ���������0����� ��P�� 0�� V�`������P���� ��L� � ��& � ����  P�  �� ��'/ ��� ��$/ � ��| ��!/ �x ��L������p ��4������h ��H������` ��@������X ��D������P �������  ��Ѝ�p���������������D ���������������'��=��F��P��Z��a��k��@-� 0�� ����3�/���� R�p@-�@��  �p@��- � �� �� ��P�⻄ � `�� ��, ���. �D� �� ������ @P�@� �� ���. � ��p����ÿ���, � ���8 � ����#���/�@ ���/��/�@-�  ������0�� P�  � ����V'8@-� @���� ���. � ��= � P� P��  | ��. � ������  P�l �  
 ��> �  P�  X ��. �  � ��= �H ��. � ��u> �  P�8 ����
4 �� P��. �  �( ��P��. � ��8����ç�þ�������������� R��A-�@��p�� `��P��  �80��  ���A�������� �� ��P��U� ����  P�`� U����� ������H �� ���������@-� ��& ���: �  P� ����N�À P�  P@-�  `@�� ����h. � ���> �4�/� �����2�À P�  P@-�  `@�� ����Z. � ���> �  ��4�/� �����i�À P�  Pp@-� P�P��M�`��  ` �� ��0��@��y� � ��� �� ����0�����Ѝ� � ��Ѝ�p���.?�À P�  P0@-� @�@�T�M�  ` �� ��0��P��a� ���$ ��' � ���� ��0��� � ��TЍ�0���.?���	���M��N-�(���=��� ��40�� ��<`��@P��D���0��8@��(p��
��< �  V� ��  
 V�&    � T�  � ��. �  �� ��. � ���� ��8��h= �0�� ��0�� 0���- �  � ���- �0�� �� ����} �  P�0�0�  0�  
| ���- �  Z�  
 ��q> �  ��  ���\ ���- � ��  �@ ���- �  Z�  
 ��d> �	 T�  * 0�� S� ��   �  ���N��Ѝ��/��ñ����������.��0�� ��������À P�  P�N-�P��p��@��;  "0�� `�� S�  0�� ���� ��< � 0��  S�    `�� U�  ���� ���
�����&� � Z�	����������	 ������/ � ��� ���  � 0�� 0����	 �ກ � ��� ���� [�p��	 ���������  �@ ��#% �<���  P� ��`@��0 ����- � ��> ���
0�� ��  ��4�/� �������	��a2��Q���N-�8C�� ����� `��K/�� ��p��m� ����; � �� ��� ��; � P��$= ���  �� ��D� � ������ ���� � Z��2�� @��  � �� �� ��/� � @�� �㰲���= � ���; � ���T���P��� @��< �P�� P�Z  ����M- � �ᄐ��z���  P�  p��2- �  ��#  � ���= � ��= �  P�  L��(- � ��  � ���= � ��9< �  Y�  
(��- � ���< �  P�  ��,- � ��	  ���- � ��= ��� Q�  
���!- � ��= � P��-  � ��= �0�� S�
  
 S�  
 S�    �!�� �� ��0���; �  � ��pa��7���P �� �����T ��  � �� P��x��- � ��  �<a����@ �� ��3� �0�� �� @��D0��  � ��	P��<���, �k ��x= ��@��T0��  S�$�  
 ��; � P� `���  0�� ��]0��0��\0��0��^0��_���@0�� 0�� ��L0������D0��  S�X ��  	  �, � ��  ����]0�� S� S` ��  
  � ��  �^0�� S�   ��
 ����0��d���h@�� ���@��< �  P�  
` ��, � ��  �0��  �� ��HP�� ��������Ú��H �á�����������	�������H�������6��V��y�Ý���F-� P��,�M�`����� �� ����p��@��V+ �  P�  
��� Y�	   ���� J�0�����  � ��2+ � P��l  �A��0��	 S�  ����}, �����0��^ ��0�� Y�1��a��:  
  � Y�
  
 Y�    �@ Y�D  
� Y�L  
  Y�7  
 P��P  �X ��$����H0�� ��  �� �� �� �� ��:��� PP�C  X�� ��$ �� a�m �=  �d�� ��h ��p0��t��� ��� a�; � PP�3  `��p ����� ��x� ���� ��% � ��t ����q� ��� ��% �#  �	 ��
�� ��0��6�/� PP� �  
  �	 ��
�� ��0��6�/� PP�x �  
  �	 ��
�� ��0��6�/� PP�
  
T ��, �  �(��� P��J���	 ��
�� ��0��6�/� ��,Ѝ�����L �����������.?����������&��D�� R��N-�@���2��8�M� ������P�� ��  ��4��  � �� ��ˁ �$ ��2�� R�   `�����+ �0�� ��0�����r����@ �� �� ��"� �0�� `��D0��r  � U�  � ��0�� �㰁 �00�� 0��: S�  S  
# S�  

 ��	�� ��0��5���  �
 ��	�� ��0��M���  P�|  ���� r�� ���XC �X ��4����H0�� �� �� �� �� �� �����  P�  � p�  
 p�  D0��  S�  
"0�� S�  ���+ �  ���+ �p ��2< �
 ��	�� ��0��G���  � p�    [�   
���� ��>  �Hq��4 �� ��X�� a�~ �]0�� S�    [�   
����$��# �  P�  
��� � `P�
  �0��@���� ��T �嵄 ���� ��W$ � ��/  ��0��` ������� 0�� E�3�/�  ��&  � ���; �0��p��^0�����^ ��0��a��  V�` ��    [�   
o���l@��^ ���9 �^ �� ��x ��^+ � ���; �  ����0���� ��  ��6�/� ���; �
 ��	�� ��0������ ��8Ѝ�����H ��(oc�����u�ï�����\%�� ���������@-�(�� @�� �  P� ��� ���� �  P�  ����·��V�� R�@-�  
 R�   ������  P�  
 P�    �"���   �	���
��� 0�� ��  P� ���+ �  �����@���) ����c�ü�� R�@-�  
 R�   ������  P�  
 P�    ����   ��������� 0�� ��  P� ����* �  �����@��) ����c�����s@-�FA � `��� ���* � @��(  �40� � ��I��.�� � ���O��.��  S����S0��.0���* �0�� 0�� S�  x0��x �� ���* �d0��0�� S�  X0��X �����* �D0��0�� S�  80��8 �����* �
 ��Q+ � @�� T�4PD� �������  ��|�����D8�Ø
��t`�í���D-�@��P�����p��  � W�a��  ��  �  �\ R�   0��c S�`� @�   
1+ �  ��`��  R� �����p�� W�����  T�  

 ��%+ �  ������@-�<0��  �� �� R�  
, ��* �  �����1�� S� ��� ��* �  �����ELF=��a���@-� `�� P��p��  � @��@��@��0�� �  
��  Q�  
0��  S�  
��� �� �� \�   ��c �  ������ ��� �����p��(`��3�� W����� ������ R��@-�`�� 2�Մ�M�P�� @��  � �� �� ��#� � U� @��   �����~ �  P�   ��F� �  P�q  ������C* ����-* �����! �  P�B\�  
 �� ��
� � P�����! � `P�  
�~ ���� P�  �!� �3 ��K � ��<  �x�� ��[� �p��! � pP�  
 ��~ �0��X��X!��  ��P� �  � ��~ �D��<!��  ��I� �8��! � pP�  
 ��~ � �� ��  ��?� ���! � pP�  
 ��~ � �� ��  ��5� �� ��! � pP�  
 ��v~ � �����  ��+� � ��`��o~ ���� P�  �!� �3 �� � ��g~ �� P� �!��3 ����� ��L���  P�  
 ��]��� @��  �x ���) � ����l ���) ���d ���) �4�/�\ ���) � ��Ѝ�����H �Ï�Ô���������	�����	���������	��!��'��0��6��?��F��l�Í�ñ���@-� @��`��p����� PP�   
���� ����4�/�  U� @��   
���� ������ R��F-� ����`��P�  
 R� P�  P�� 0��- S�  
 �� P��  P�  
 �� ��g � @��  ��0�� @�� ������  P�@�2  
  U�   
0��p S�P� p�P�     � �����  R���  
��
 ��~ ���� ��0�� �� \� l�   
k~ ���
 ����� P��2�� W�p������@��  � ������ @����4 ��d) � ��I� ����� @�� �� �� @T�@�Z) � ������H �������� R�@-� 0��  � �� ��
 �� � 0�� ��  c���� P��@-�P��@��� ��,  ��� �� �� � `�� �����G � pP� �  
 �� 0��  S�  
: S� �	   �� �� �� ���~ �0@� S� P��  �h ��) � ��  �P����T �� ��) � T�  � ���� ��b �  P�  
, ��) �  ���  ��) �  ��������=��Y�Ç�î�������� ���� ����� ����  ����� B��N-�@��p�M� R��-  � ~��P~��x~�Ø~�����  �  P㸲�  
 �� ��~ � ����� ���  � �� �� �����~ � �����r  � P��  � �� �� �����~ �P�� ���  � �� �� ��~ � �� ��P�� ��� ��~ � ���  �w' �  �  U�  ��( � ��}  �l�� �� ��~ � �� p�� ��eG �  P� ��  �� �����( �����l �� 0��  S�`�	  
: S����� �� �� ��l ��w~ � `P�  
����� �� �����8G ����  P��p�
  ,���h��  �����
 ���| ����  P�  
L��
��( ����� ����0��4�����@��( �  �$���� ��0��( � ����Io �  P�� �0�� �  
�k �  P�  �� ��� ��0��n( �  � ��n � �P�  ���� ��f( �  �  Y�
 Y ��	��1
��m �
 P� ���  
 ����0�� �� `��V( �<k ����:k �t0��`@��	��l �� ���M( �	 ��`�� ��|� ���T ��! �  ��pЍ������	��  ���	����N��t��/��G��N�Ã�ó��������%��(+��H ��;��J���� R��D-�@��P��  ��& �  ��� �� ���} � �� p�� ���F � �P�  �� ��� ��( � ��.  � �� 0��  S�`�
  
: S�  
� ���' ����� �� �� �� ���} � `�� T�
 ����t@�@��n �  P�� �0�\ �  
Ck �  P�  �� ��D ��0���' �  � ��,n � @P�  
( ���' ��j ������j � ������M��s�á�������ã���/��/��/��/�0��  �� ��  �� ���/�(��0�� �� P�0�2( �3  �#�0 0�/�(��0�� ���/�(���@-� `�� @��  �@| �P��(0��T%�@�� p�� ��9| ���  W� ��  | �  P�   ������P�� ��0�� T����:  ������(��7@-� ��' �1�� 0�� S�  � S�	  * S�  
 S�	    �S�    �� ��  �� ��   �� ��' �� �� P��' ��@��)  �� ���� ��' �  U�  
 ��0��0��  
�!�� ��' �  � ��' ������0��	  
 ��0��,Š� ��ˌ�!�� �����u' �  �h ��r' � 0���\ �  �T �T �j' �P��(@��H0��0�� U����:>��� �����4 ��< ��7 ��>V��8��E ��W ��c ��n �� �È �Ñ �Ëd��(��@-�0@�� ��0�� S�������(��� ��� �f| �0��0��0�����(��@-�  ��@����} � �� 0��M S�  
  �K S�    �k S�  
m S�   �� �� �� ��  T� ��0� 0����4��$���N-� ��A�M�x��  Q��M��� ��  ��� � @P��  
�{ ��? � @� R��  �P���� �� @�� ��.| �,��' ��  �Am�� ��`��P&������� �P���  
��D �� 0��@ S�  *�� ����D �����:��D�� 0��( S� ���  �  ����  ���  ���)���& �  ���� P��0��D0��ʍ� ����D ��?{ ��� ��  P��\�D0�0�  
:��D ��4{ �d�� ��  P���\�D0�0�   
ʍ�D ��){ �<�� ��  P�  ��P��D0��0��D0��	  �:��D ��{ �  P�  ���@P��D0��0��D0��ʍ���� ��D ��{ �  P��D0�0�D0�������  V�(��� ���0���8P��4���,���N  
pf� W���K  �
�� ���� ��z �A-�� ��
P��p��0�G�6  � ��������0���Р�������� `��1  
ʍ��!��0���� L� S�
  �    R�  �ء�������� [�#  �    Z�   �С��
 ���� Q�  �	   P�  �ء�������� Q�  �  
 P�  �z����p�� ��z �  P�   ����z �  P�  
P��X1�� 0�� U�����H1�� 0�� U�?  �  �l��S& �  ����DP��  �X��M& �1��  ��1�� ��#  � 0��  S�	 S  

 S�  
 S�  
, S�  P�� U�  *���� U�*��:  ��@�� 0��' S�  ��P��� ��0& ����  �� ��J{ �  ��(�㼖 � ��  �� ��%& �   �t���  ��HЍ�ڍ�����`��ʍ�)��D`�� ��z � pP�+��&��������0���Z��P��t ���`��� N����`��8������	& � ��������� ��(�õ �ý ��� ��!��A!��l!���e�â!�è!�î!�ßd�ô!���!���!��0�� "����P"��k"���N-��M� @������� �� ��E���z �0�� ����  
  R�   Z�  �����% �  �������% ��0����� ��1�� � 0��(�  
 ���!��& � �P�%  
�0��4p����  �� ��1��t`��TP�� q��$a��(Q���~ � �� ��l���~ � ��0�� ��X��$��+��4���~ � ��0�� ��8��$��+��4���~ �  �� �� ��E?�� ��  �`��P�� ��0��d�����T��k��[��% ��� ��) �{��'{�� ��� ���H �  W� ���  
��+g�
0�� �����������o��% �[E�`��P��k��;��#;��  S�  
�� ��c�  ��
0��������\���_��u% �P��
 ��' �%5��(  
4���Ԑ��� ��4��t���Tp����� ���$���(q��~ � ����~ �	 ����  ��~ � ��
 �����~ � �� �����~ �$�����!�� ���(��� 1��������M% �  �� �� ��E?��_ �  ���E% �0���� ��4����*& �  ��   ��  �K_��l��`�� Q�� ��a��4p��$q��d~ � ��T��y � �P�  H2����� Z�  �0��8��
 ����� ��1��$Q��P��(q�� a��Ay �
 ���� ��=y ���	 ��I~ �	 ����  � ����� ��P��2y �:  � �����[y � �P�  �1��(�� R�A�P�/  �0��`���� ��$Q��1��P��(q�� A��y ��� ��(~ � ��	��5 �  � ��l��?y � �P����
 ��\��:y � �P����
 ��L��5y �  P�A�P�  8�� �� ��P���x �/��T0�� ��/����� �� ��(1��~ � ��4 ����~ �  �� ��E?�� ��f �0��8�� S� P��   ����y �  P�  
 ����y �  P�	  
 ����y �  P�  
 ����y �  P�  @��x�� ���} � �� ��r5 � e�ލ�����"���"���"���"�������"��	#��)#��J#��P#��2r��U#��i#��7%��  �#��a�Ô#��M�Á�à#��'�å#�ì#���N-�8�M� ��0���5�� ���%�� 0�� S���  � S�  * S��  
 S��    �S��  �  �E��4���  ����`��	 ��} � 0��|�� ��0��(P��x �0�� ��� ��� ��x��C#�T��b ��������0p�� ��|x �0��8�� ��C#��b ��������0p�� ��rx �0���� ��C#��b ��������0p�� ��hx �0����� ��C#��b ��������0p�� ��^x �0����� ��C#��b ��������0p�� ��Tx ���� 0��	 ��������L,�0��� ����� �������� ����������0p������ �00�� S�   ��xG�P��` �:x ����(��� 0��$���	 ��N,�,��勴���� ������ኤ�� ��� ���0p��$��媻��,��労�����(���0��������� ��� �00�� S�]   �����` �x ����(��� 0��$���	 ��N,�,��勴���� ������ኤ�� ��� ���0p��$��媻��,��労�����(���0��������� ��� �00�� S�;   ��H��` ��w ����(���	 ��$���0���N,�,��� ��勴�� 0������ �છ���� ���$��� ���0p�媻�� ��剤�����,������(������o �00�� S�   �����` ��w �0��,���$�� ��C%�( �� 0��Ġ���ˌ�$����4��0p��$��� ��  ��,��(0������  �d��@��# �\��  �q���  P�@��  ��� Z�6  ����8�� ���w � @P�  ��� ������ PP�  �� @��# �o  � `���� ��@��r V� �� ��f� `�My � �� �� �����`  �0�� S�  ���
 ��0�� ��oy �0��0 �� ���Ϡ� R� ��� ��  \�  
 ����c# �`����� 
� ���  � ��� ��� `��@�����X���Z �  P� P�:  ���� `��p��
`��p��_Z � Y�  � 0� P��  ����  ��0��  U�  
 ��0���# � ��0��  P�  ���B��  T�  
� ��  � u�  � ��P��2# �@��  � U�  � ��,# �  � U� P�P	  U�  
 W�����   V������ �� P������ Y����`��p������U �  U��� ��8Ѝ��������(��2r��M�Á��7%�à#��v��'��q;�ù#�Ë���#���#���#��$��$��4$��� ��]$��u$�Æ$�ä$��02���N-� �R�`��$2���� ��0�� 0�� 0�  �0� 0���� ��P��������`  �  U�  @�� ���# T�  
  Y�  
 T�
 T ����p�@��� ��p�@���b  �	 T�  T\  
 T�Z  

 T�p�@�Y  U  �pr� p�3�q� ��3@��  
@�� T�
 T    [� @�����p��  ���� �F  �  W�  
  T�	 T @��p�>  
;  �  \�@��  
	 T�  T p��4  
4  � T� p�p� T�
 T-  @P�\ T�    W�  
���
 \�����@��p��  ����� �� @�   �  P�  
 �����  [�P�� �� ����0�� �� ��� S���:  U�  
  [�  
  R� 0� 0����  Z�  �   ��,��{ � ������p��@������� ��P������� ��(���$���F-�`y����M� @��P��  ��  R�C  
  Q�<  
0�� �� c� U�P�!,)�� �� ��  ��uw � �� 0��P��P�� U�  :0��  ��P`��P@�� S�  ���� ��� �y{ � ��v �  �� �� ���Y �8�������<" �8�� ��  R�# 
 ��  Q�  
�$��&��  R� 0��  S����," �h8���� ��6� � PQ�p�   �h��"" �d�� " � �P`��X�� ��N{ � ��L�� ��gw � �P�   ��8��cv � PP�0��2�� 
�7�� ��
��
P�� ���v ���� ��8{ � ��}v � �� �� ��Y �
 ��
��
 ��
0������ � ����� ��Ew � �P�.  @���� ��v ��� ��=v � PP� ���	  
 ����6v � PP�  H7����  Q�� 
 ���u � �l�� ��*v � PP�7�����
 ��P��#v � PP�  �6�� ��  R� �4�� 
k � ����oS �
P�� � ���� ��w �  P�A   ������ PP� ���~ 
�6�� 0�� S����  
 C� R������  � S�  �����! �6�� 0�� S�  
0C� S�  ���� ���u � `P��  
��� ���u � `P��  
 ��|���u � `P�  p�� ���z � ����S2 � ���  Y�  
P ��L��z �e ���@��! �	P��P ����B � ��(��	 ���v � PP�  	 ���� ��Cw �P��P�� 0�� �� 0�����k! � @��  T� ����  
T5��0�� T� ����� P��% � �� ������  � ���� ��v � PP�P�b  0��S�[  � ���5����p���0���P�����P��H! ���x��E! �0����� ��h��h%������0��pz ������ ����H��Uv 멕��8�� ��8%������Ѝ�cz ��� ������Iv �p�� ��[z � ��u � �� �� ��X �����v � 8�����(���#<��4��"4���$�� S�  @p�����! � ��u �  P�
  
�ğ� ���� ��0��p�����ğ��P������ �  �� �� ��  ����  � ���� ���0������h���  �d���  �P ��\��%z � P�� ��P�� ��=v � �P�  dc��p��  W�  P ��,��z �P���  �@�������/u � pP�J  ,3�����@�����  ������  �������0�� ����  
 W� ��   R�L  �43�� 0�� S�
  
 S�  
0C� S�  ��2�� ���������� P����`������0�� ����  
  R� ��   R�1  ��2�� 0�� S�  
n�� S�`��e����  
0C� S�  �@2�� ��0������� P��  U�P`��� P�Q  ������  � ��9  � ������ @P�  @��P ��y �P��k  �0�� �� Z�0��	   R�  �  S�  
 P��[�  P ����?  � P��[�   
�"�� ����y � ����  ��q���  P�  �� �� ��k��� PP�
  
�� ��D��`��a  �<��P �� P�� ��y �>  ���$��X  �P �� ��  �d1�� 0�� S�3  
 S�  
0C� S�.  ��0�� ��P`����U��� pP�  
�����B  � �����  �����<  ��� ��P��ky �  � ���� ��u � `P�  P@����P�� ��_y � ��t � �� �� ��W �\�� ��Vy � ��t � �� �� ��  � P��P@�� ��t �  �� �� ��W �   � P�� ���Ѝ�����(��� ���$���$���$��K�È��Ëd��%�� %��*%��/%��6%��B%�ö���J%��N%��V%��_%��"v��l%��s%����Ð%�ê%�ù#�ø%�Ë���%���#���%���%��&��%&��/&��N&��d&��w&��c��;�À&�Ó&������ � @  �@@B V'�&�ù&���	���&���&���&��
'��!'��('��v��'��x'�å'��@'�ý'��X[���'���'���'��b'�Ç'��(��
(�� R�s@-�@�� ��*  ��� �� ��u � P�� ����g> � `P� �  
 �� 0��  S�@�  
: S�  
p �� � ��  � �� �� �� ��{u �0@� @�� S�  �@ �� ��� ��4 �� � ����ck �  P�  
 �� �  ��|����(��)��4)��b)�Ê)����� R��D-�@��  �� �� �  ��0  ��� �� ��p��Uu � `�� ����*> � �P� �  
 �� 0��  S�P�  
: S�  
| ��` � ��  � �� �� �� ��>u � P��@����P ��h �
 �����j �  P�  
0�� �� ��, ��^ �@��$ ��[ � T����Kg �����)��=��s���)���)��*�� R��D-�@��P��� �� @��/  ��� �� ��u � �� p�� ���= � �P� �  
 �� 0��  S�`�  
: S�  
� ��@��! �  � �� �� �� �� u � `��
 ����j �  P�  
�� ��0��@ ��$ �@��  � T� �, ��j �  P� @��  
 �� � ������4*��=��s��g*�á�Ð*�� R��F-�d���M�`��@��	  ��� �� ���t � p��\B �F � PP�  
0��� � ��F  � ����= � �P��  
 �� 0��  S�P�
  
: S�  
� ��� ����� ���� �� ��t � P��
 ����\j � �P�  
�� ��0�� ��� ����� �� ��
��t � V�
 � ���   ��
�� ��t �  ��	�� ��2j � p� `��   ��0����T �� P��� �����@�� ��@ �� � ��8�� ���w ���, �� �  ��Ѝ�����*���*��=��s���*��'+��Q+�� ����@-�4���4@�� ��0��0��@l�$�� ��  ������ ����� ����|�ì�ë���  ��* R��/ �� �� ��bt �@-�  ��@��* R�   �� �� ��Yt � T� ��� T�  ��� T�  �  �  ��� �� ��Kt �A�� 0��������N-�@�����`�� p���r 봱��Q�� ���a  � ���r �  P�\    ���r �  Z�X    V�P��,   ������ @��	 ������ p�� ���r � `�� ���r ��� P�  �1 �! ��r � U��(  �ب������������������ p�  �3����  P� �����������  P�  �� ������  P�  �� ������  �������� ��������� @��	 ����� U��  �l���|��È��Ø��è��ø���  ������  T�  � �����  T� �����  T�  �� ������  T�  �� ������  T�  �� ������  T�  �� ������P�� U�
 �� ������ �� �  ������|�����-�� R�@-�@��  
@�� ���  �� � �� 0�� R��  �X���p���p���P���P���p���P��� ��  � �� 0�� ����k���  � ��� �  �� p�  �3���.��`0 �@ S�  �/0 �? S�@ ��/� 0�� ��   � ����0��  Q����R3�� ��? ��/�0�� �� �� ���/����0��  ��  R� � � ��/����@-�0��  �� ������������0�� �� �� ���� ���/����0�� �� �� �� ���/����@-�@@�� ��  R�  
������ �� 0��  �$ ��  R�  0��0������� ��������$0��@-�(@��  �0��, �� �  T�@D�����������8@-� P�� @������   � � ��@��  P����8���1��  ���A-�A�� `��0 ��G��, �� P�( ��F �0 �0P�����#��-���$��40��Pc�  U� ��@  �PU�~0��L0�� �;  
PU�!0��M0�� �6  
60��PU�  ��N �� 0C� ��0�(0��-  
7 ��PE�o���  U�@0��O0�� �, ��$  
PU�80��- ��P �� 0C� �-0��  
90��PU�# ��Q ��	 �$0��  
PU�N0��R0��
 �  
PU�1 ��S �� �  
 U�T0��0� � �" �~�U �  �X�V �W�\@��p�� 0��  ��`�� P��I ��I ��J0��0��H0��X0��K0��HP��=���0��- ��0�� ��H ��H��IP��H ���A��������p@-�L@�� 0�� P��I �� ��J0��N0��H ��" ��K0��I ��LP��$���-0��NP��M0�� 0�� ��L0��p@��m��������p@-�L@�� 0�� P��I �� ��J0��Y0��H ��" ��K0��I ��LP�����-0��NP��M0�� 0�� ��L0��p@��U���������@-�C�M��M� P��B��B����0��$4��; � @P�`�  
  �@���q �B.���� �� ��\: � ��p���� 0P� ��`�� ������  �,�� @��>9 � ��d �� �B��k�� ��?9 �  ��L��r9 � ����E����� ��4 �� � ��,�� ���u ���  ��t � ��4Ѝ�ۍ������7�è��Þ.��J����@-�" �  P�    �����@��" ��N-���(�M�@��`�� �  P�T�  
 �� ��Pr � P�� T�p���  � �� �� ��Hr � T� P���   �� ��
 ��Ar � @P��  
 T�  
����i �P�r �@��2 �P�r �� � P����  ��x��p � `P�  �� ��d��W � �����  ��� ��L�� `��O �D3��# ����� ���$ ��4#��P��(`�� ��(#��,`��  �� ��- ��������3��4 ��0 ��� � P�  
 P����t  �� �p���� �^  
� �p �� ��� �Y  
 `@��`�
 V�  ���   �u��� �p���� �L  
 �I� ������K�	��� {�
���4  � �p0��� �@  
 0�� �p���� �;  
� � 0��p ��� �6  
	������Y#��	 ��? �  �� P�.   0C�_ ���0� �K�	�����{���  � �p0��� �"  
D Z�   �� 0��Q��� 0��	  �S Z�  �!��H���0 �� ��0�� Q�0��0 �%����K� [�����y �p ��� �	  
Y3��	���?�	� ���	 P�  o �p �� P�  
������)��� ������
`��
  �S Z�   �����R���  � ������B Z�=  
��������� `�� ���O ����  P�   
Q ����mq �d Z������� ����P����� ��� �� � �����
 ���t �
��� �� � u㸠��   0�� �� 0��`�� �  � ���� `�� � P�� T�  
�� �� �P�Gq �p��H1 �P�Cq �$ � P���� ��(Ѝ�����@��%��� 0��D ��`B������	��  ���.���.���.��=/�����ܪ�����Þ.��J����H ��|/�á/�ÿ/���F-� `����M� p��P�� @��F  � �����3.��!>��_0 �  P�e  � @� P� �-  ꘴�Ø��Ø���,���,���,���д��д��д��0���!��4#��
���
 T�
@�!
 ��mp �43��0C�
��� Z�  �  �`���`d��p �1~�� ��0������ `��> � �������� ����� ��jt ���� �� �0��4  �����0�� 0��  S�  `��d�� ��ǌ �  Q�  . �� �
P����� �0�� 0��  S�p���  
	 �� � Y�  
  �  Y�  
  �
 Y�  
 Y�  
 ���P0�� ��T0�� R�  
� �  P�	  ���?�� Z����:0��  ��
0c�  ��  S����  ���ߍ������/�� ����|��T$��8@-� ��@��P�� �  P�  
 0��1 S� �   
  ��0�� T� @�  ��   �� �� ���p � @��p �� P��� � ��h��� @��j �P��  P�   
l ����p �d U���� t�  0 ��� � ��8�����  ��� �0��  �� @��8���T0��|��_0�Ã0�á/��H �� R��D-�`��@��  ��D��d � �� �� ��p �h0�� �� �� p��p�� ��}p ���  �� ���  ��/i � J��� �� P��, ��0�� � V�  
 �� �� ��kp � P��  ������ ���1�� R�@-�  � �� �� ��_p �0��  ��0�� �� �� �  ����� ���1�� R��N-�P��`��V  � �� �� ��Lp � U� ��Q  
 �� �� ��Ep � U�  ��L  
 �� �� ��>p � U� �� @��  
 �� �� ��6p � ���P�� ������� �  P�"    [� Z  �J�� ��	 ��W �  Y� �*  �� ����� ��P � ��0��  � �� �� �� S����:� ��p��1 �`��  �  �� R�  
? ����� �  P�  

 ��� � ��  �p��`��  ����0��L �� V����:  T���� @d� Pe�@���������1��0�� �� �� @��������2��a2��92��b2��m2��  �E R�p@-�`��  �p@��� �  ���� � PP�0  � �� �� ���o � �� �� @�� ���o � P�	   U�   0������ U�  �0������ 0������ U�   �� 0��  ���0C�  S����
���� U�   �� 0��  ���0C�  S����
���� �� 0��  ���0C�  S����
���� ��p��� R��G-�P��  
�G�� ���  ��m � @P�  � �� �� ��o �`�� �� �� p�� ��� ��o � �� �� ��� �� P��o �  P�p���  D �� � ������ T� 0� 0�  
 T�0� 0��0� 0� P�p������������ �ß2�� R��D-����  
Ѝ��D��O ���  ��8 � @P�P��J  � �� �� ��`��ho �Q���� �� p��p�� ��ao � P���� ��P�� ��[o �$  � T�
    �� ��� R�  
0����� ��P�� ���} �  � T�  � ����� R�  
��0�� ��  �  �� ��� R�  
� ����0�� ���P��h �
  �`��p��P�� P���� T� P�   P��H ��  �D0�� T�@ �� �<��� V�80����4 ��0�Q � ��Ѝ����� �ð2���2��&3��e3��\3��a3��a2��Y[��j3���G-�@�� B�P�� R�  ��G��� �  ����� � `P� ������ �� �� ��o �h0�� �� �� ��� ��� ���n � T� p�� �   �� �� ���n �	���  � V� p�  
 V�p� p���� @�  P�������� �� S��F-�(���p��  
� �>  �a����0 ��    ���� � PP� ��4  � ��	�� ���n � @��@����� ��� � U� �� �  
 U��� �� � �� � ��E- �  P�  
 P�
  �0�� 0��- S�    W����
  P� 0e0�@������h`���� �� ��n �0�� S�	  
 U�  �  
 U� �  �  W�@���������0��  ��0 ������ �Ë3��!v�Ò3�Ø3�Þ3���6�����@-� �� 0�� ��0�����������@-� �� 0����0���������N-��p������0�� R����`�� P��@��  �Ѝ��N��S ���    ����: � @P� ��  � ��	�� ��kn � `�� [�`��  
 ��	�� ��cn � P���� �㤉 ��� ��0��  �� ��d&�Xg �0�� ��  ��@�� P��`��Ѝ����� �À���A-� P��  ��`��p����� V� @��  
 ���A�� � �� ��
 ���_��=n � �  � �  P�d ��  
  ������n � ����� P����:  ������ R�s@-�  ��  � �� ��
 ��&n �; � @P�P�Q  
 0��0���? � PP�  
4��J �I  ���(��F �o�� ��C �l����Q��? �p���l��\8����,,��\������ ������5 ���� ��2 ���� ��/ �0 ����������0�� ��R"���& �<���0��� ��  Q� ���� �����`�孈 � �� �᪈ � �� �� �� �@0�� S��	  
 S�x�  
 S�p�  
l �� S�h���d �� ���\ ����� � ��|���6���6���6���6��7��7��$7��qj�Á���67��H7��K7��O7��b7��z7�À7�Æ7�Ð7�Ö7�à7�ï7���N-� P��`�� R���  ������������È��������������� ��|��)l � @P��  ��
 �� ��m �); �  P��  
`��~? ��  � ��D��l � `P��  
 ��; ��  � ��(��l � @P�;  ��
 �� ��m ���
 �� p�� ��m ���
 �� P�� ��m � @�� ��; � �P�  
 ������k � pP�`�d�  
 �����k �`��  P�  
��� �p��0�� S�  ����@��@��� �  T�  |����@��@��� �
 ���� ��0���9 � `P�T� `�P�� �  � ��D���k � @P�:  ��
 �� ��Km ��� �� ��� ��Fm ��� �� ��� ��Am ��� �� P�� ��<m � p��	 ���: �  P� ��h  
���	�� ��0��` ����`d��?� V�`�!��
0��	 �� ������� ��  V� @�� p���������<   U����� ��������`T�`���X��;  � ��P��k � @P�<  ��
 �� ��m ��� �� ��� ��m ��� �� ��� ��m ��� �� P�� ���l � p��	 ��: � �P�)  
� ��	�� ��0��! �`d��?� V�`�!��
0��	 �� ������  V� @�� p������  
� ���� �� `��	  � U�����| ��`T�`���p0�� T�l �� � �  ���`��X ��� �   �`�� �������7���7��J#��c��P#���7�� 8��8��38��I8��^8��c8�Ò8���"�é8���8���$�æ8���7�� R��@-� P��@��#  
 R�G   ��,��-k � `P�B  ��
 �� ��l �-: ���
 �� p�� ��l ���
 �� P�� ��l ��� @�� �� ��8 � `P�� �)  ��� ��� ��� ��(  ��� ��k � P�  
 �� ��l �: ��8 � `P� �  � �� � �� � �� � �� �| ��  �x�� ���j � P�	  
 �� ��ol ��9 ��8 � `P�P �P �� �  ���`��@ �� � ������&��<9���8��9��g9��Q:��l9�Â9�Ó9���9��:��f:�Ã:��l:���7���M���8@-�4@�����  T�,@�� ��;��  �  �_��  ���� ��0��,� � �� �8@��Ѝ��/�@-�L ������$!�� �� ������F-��0�� p��@�� P�0�� 0��$0��$0��  S�P���   
  �
�� ��i� ����P��?`�0��  �	 S� ��`�����P��`��@ V����P��U�  
���`�������3 �0���0��0��?0��0���� �� �� ���0�� ��� � ��� p�� �� ���0������}�� �M��N-�(�M�p��H���l�� `��p@��  Q� ��X��� ��$���\P��d���E  ����-� ��� �� �᱇ ���� ����%� ��� �� �ᩇ � w�����  P���X���\P����� ��d���`f� �� �� ��$���� �� ��u���T0��	��
��J�  �� � `�� `��$ ��� �P����� ��<  �`F� p��p��	��$p�� ���� �	�� �� ��}� �`�� ����� ��� �� ��u� �����&  � w�0��  ��0�� ���# �0�� ��� �� ��? �� ��  P���X���\P���� ��d���`f� �� �� ��$����� �� ��5���h0��0C�0`�$0��`�� `��  �`@� p��p��$p��(Ѝ��N��Ѝ��/�8@-�@�� �� ��uk � P���8 � �P�  0 �� �  ��8��� ��0�� �� ���� �� P�  �  �8���9<�� ��@-� ��^k ��8 �  P�   �� �  ����� ��0����  ����9<��p@-� P�� �� �� ��Kk � `���8 � @P�X � @�  
0�� �� �� ������ 0��0�� P�� ��= � @P�  
 ��e �  � U� @� @� ��p���9<�ó6��p@-� 0��P�� @���� �� 0�� ��0��0��pj �  ���� ��p@��kj ��L-��M�@��P����p��Hb�����  P�  @D� T��  �������H���P���o��   �s�� ��������2�����  �� B��ʿ������_���@�� 0��  �w������{������  ��ߍ�����0@-��M�@��P�� ���� 0�� ����� �������D ��H0���� ��)��� �������l ��p0���� ��Q��� ������ ��0���� ��y@�� @������� � ��  �$ ��  R�  
(��  Q�  
΁�	������0��� ���� ������� �L ��  R�  
P��  Q�  
΁�1������0�� ���� ������� �t ��  R�  
x��  Q�  
΁�Y������0��d ���� ������� � ��  R�  
���  Q�  
΁�������0��, ���� ������� � ��Ѝ�0���d��X<�á<���<��=��L=���M�@-����0@�� �� ��0�� ���� �� ��B���	 �� ��0���� ��  ��;���$�� �� ���i � ��(�� ��i �@��Ѝ��/��N-��M��P�� @�����`��( �� �� ��,0��i � ����p��)��������@�� �� �� �� ���� �� �����  [� ���  
,0�� �� �� ��Mj ��� ��� �� �� �� ��,�� ��
��  � ����� �� �� �� ��K�� ���������� ���|0��8���P��90��8@���p�� �� �� @��	@��4@���@�� �� �� ��	 ���� ��)���
 [�  
,���
��
 �� ��j ��� ��� �� �� �� ��,�� ��
��  � ����� �� �� �� ��K�� ��������� ���|0��`���`@��a0��P���p�� �� �� @��4@��@��0@�� ���@�� �� ����4 �� ������
 [�  
,���
��
 �� ���i ��� ��� �� �� �� ��,�� ��
��  � ����� �� �� �� ��K�� ��������� P��|0��P��8���0��@��P���ؐ�� p�� �� ��� �� �� ���� ��0 ����������P��0��0��x��� �� ����� �� �� ��00�� �� �� ������� �� ���h �H���s��Up�� ������q��`p�����U��������� �� �� �� �����p���w�� ���������� �� �� �� ��������{��p�� ����������oo��`�� �� �� �� ������������� ��`��`�� �� �� �� ������ ��܍�����p@-��M�@��,�� �� `�� ��P��h � �����  P�  � V�  � ���0������ ������� PP�	  , �� �0��p �� ���� ��h��� ��   �  ��܍�p���=�� R� Rp@-�@�� `�`�P��   ��X���g �  P�   ����p@������ ��8���g �  P�  �p�� ����p@��G��� ��j � ��h � ��p���=�Ü=�ß=�ÿ=���F-�p��0��|�M� ������ 0��r S�  
w S�  
i S�   � P��  � ��  P�  
 ��
 ��i �P�� @��  �� �� ��yl � ����$ �j  �P��0�� ��
 �� `��z`V�`�0f���	i �0f�1�� 0��k S� @��  
  �b S�  
f S��    �t S�  
u S�  
r S��    �0f� Z� ��  
�  �0f� Z���  
�  �0f� Z���  
�  � Z���  
�  � Z���  
�  �0f� Z�  	���0f� �� �����h � ��� ��Z6 ��� ��`���  Z�'  �"��
0��(��  ��  Q�  
0�� S�������  U���� �����b��2��p�������0�� p��� ��  U���"��0��
 �� � ���� ��l �
 ����# �d��� � ��  � Z�  ,"�� 0��(��  �� Q�  
0�� S������  U� ��������b���1��p������������ Z�  �!�� 0��(��  �� Q�  
0�� S�������  U� ��������b��1��p����������� Z�  t!�� 0��(��  �� Q�  
0�� S����T��  U� ��������b��@1��p��@��X������� Z�)   �� �� ��[h �1�� �� `��( �� 0�� R�  
�� Q����� ��;�� ������0��r��  U�� ��d�����`��0�� �� �� `��o ����  U� ��0��
 ���� � ���p��`�����	 Z���h �� 0��(��  ��	 Q�  
0�� S����H��  U� ��������b��40��p��4��T ���c�����H ��J �  ��|Ѝ������>���������>���>���>���"��?��^8�Î=��2?��[?�Ê?�õ?���?���7�� ��  ���/�  �� ��  �����/� ���������� 0��  ��  ���� 0��0���/� 0��  S�  � ��/�@-� 0��8 ��  ����@�� T�  	��� \���  ����� R� �����  �����4��@-�  P�  
�0�� Q�  �1 ��30�5  : ��0�� S�L �  
H��� S�D �� ����	0��8 �� ���� �  � Q����  
 0�� S� �����  �����+C��(C��$C��0C��@-�0��@��  T� 0�  �    � S�
  0�� ��p��@�� ��r ��	k ���\ ��
 �  ��� 0�� ��r ��8�� S����,0���� �������  ��� ��
 ��� ��
 ����4��2r��bC��lC��1�� ��  S�!/�4�  
�4��6��  S�"*� �  
;��#;��  S�"%����j �wC��{C��C�ÃC��0@-�P���M�@��  T�  
0���� Q�p �  
l �� Q�h ��  �TP��@��	0�� ��T����� ���j ���D ��a
 � ���� ��e �  �( ����Y
 �@�����Ѝ�0���4��+C��(C��$C�ÆC��&���D-����`�� @��$ ��
 ��K��� pP�  
 ��
�� ��5���0��0��0��&  ��0�� �� T�  �� ��R��� p��P��   � ��0�� S�    S�  � ��T � ������  � �������0��  W�0��0��	  
 ��0�� R�  �L0�� �� �� �����   �V���  ������ P��
 U���� �������0��0��0��J���  ������4�ÎC��p@-� @�� `�� P��  ����� ��� �@�� P�� T� �����p���8@-� P��P@�� ������ ������ �� �0�� U�   ������  P� � 0� 0�0��h���   �"���  ��8���4��@-�  ��@���f �  �� 0��M S�  
  �G S�  
K S���  �k S�  
m S�  
g S��� �� �� �� ��  ������@-�@��P��  �����p��  �� �� `�� ��?e �  P�0� �  �0�  
 �� ����5e �  P�0� �  �0�	  
 �� ����+e �  P�  0�� ��  ��0��0�� ��d �� 0��0�� �    ���L ��  �H ���� � ��  ���  ��f �  U�  �� �0�  � 0�����+C��$C��(C��H�÷C���C���F-����1�� p��P��@�� `��  � 0�� 0�� `�����  � ��� ���d �  P�P  
 0��0�� 0�� ��� 0����0�� Y���� `��1�� V����`�� 0�� �� 0�� 0�� ��p&��� 0��0�����  P�
   0�� ����, Q�  ��  0��  S�  � ��q � ��)  ���>f � 0�� `��  V� p��  
�� ��e ����� ����A���  P�  ��  0�� S�d�  
` �� S�\��� ��T ��S �����wp����B���  P�  �� ��� p� �  ( ��G � �����������4���C��D��+C��$C��(C��6D��KD�� P�0��0@-�P���M�P �  
L�� P�H �� �D�� ��ai � ��{< �@��
p�  ��  ��  ��� ��$ � ��Ѝ�0���+C��(C��$C��^D��cD��0���N-� s�@�� P��0� �0c  ��0�0�� R��� ��z  ����� Q�  �0�� S���  
�!�� S�����	 ��0�����j  � Q�  ������� �e  � �� 0��0"� ��	�����  P�]  0�� ��  ��,���  \� `�'  `�� ����� �  Q�  
0�� S�H�  
D!�� S�@���	 ��0��<��C  ��� ��� �  Q�2  �0�� ��� ��� p�����  � �� R�  �  
 ��p�� Z�������:`�� �� V�����0�� S��  
� �� S����	 ��0�� ��  � 0�� `��p��  ����
��� Z�  
���
0�� V�`�����: ���� P������� �� R�  
0�� S�4�  
0 �� S�,���	 ��0��0 �� � ��   �  ������yD��+C��$C��(C�áD���D���D��NE��E���N-�(�M� pQ� 0��:�� 0� 0�� P��0�� �� 0��0���c � @P�4��  
04���e� `��
  � ���c ���
 ��  Z�   ���c �  P�  
 `���3�� V�����  �@��;�������� ���c � ��	��8���p��  P� �0� �0� � �  �� ��  �$@�� 0��- S�@�$@� ��  
 ��$��;���
P� ��� �1h�59  :$ �� 0��@ S� ��  (�� �� !�-��� ���$p�� 0��( S�`� p�  p��)��$p�� ��c �  P�$ ���*  
`g� `�� V���%  
 ��$ �� �����$ ��wc �  P�$0� 0� �0�0� �$0�$@�� ��, Q�   y��  
@��$@��  �; Q�  Q  
��� �D  �( ��  �� ��, �  �� PP�  l��� �:  � ���c �0��  W�( �����0����� ��  
�� F�c � 0��  �
0��	 �� ��h �0��0�� ��0��`�� 0��0F����0�� ���� s�0� � ����� �P�  0�� �� ���� �� ����� ��0��s0��0��  T�  
 0��  S�  
; S�s�� Z�`��p��   �����A  �0��  S�  0�� S�\�  
X!�� S�T���0��	 ��H�� �1  �  T�  
 ��; Q�    W�@�    �  Q�    W�  
 @��  ��� �  W� 0� 0�  � ��� � @P�  � �� �  � �� ��c �  ��`�� �� ��N��� ��L���P�� `��  �S����� ��P�����  P�  
 ��W��� ��  � `��0�� �� U����0��  �� @��(Ѝ�����
�� ��D ��h �����G��4��T�ÅE�åE���E�Ñ#���E��F��EF��TF��+C��$C��(C��dF�ÈF�øF��@-�0��@��  �� #� �����  P�0� �0� 0����8@-�@0�� @�� P��  ���� ����� ��� �@�� P��0�� �� T���� ���  ��8���4��0��  ��@-� ��( �����@������4���N-�lE��(�M�(R��  U�    ������ �������� ����c ���,��( ��c ��� �� ��c �0��(2���� � P���� � @���� � 0��0�� P�  
 �� ��)b �  U����  
 ��zb � P�������
  �  T�  ���� �  � ��ob �P�  :������ �  �|��,2��  S�  
����9b �  P� P��  
T4��P�� `�� p��  ���� �� �`�� p��,4�� ��  �� V����  ��,"��������X  ���' �� 0������  P�Z  0��  ��= R� �3  ' �� �� ��0��0��i���  P�Z  ���,��	 ��)b �  P� ���i0� ��0�  	 ��+b ����  Z��  
t��'0��  �� p��  ��� Q�  	�� Q�  
 p��l�� W�����  � S�\�  
X�� S�T�� �P�� �"  �H�� �  � �� ��b �  ��0��	�� J� ���	 �� ��'���0�����0��0��a �0�� ������J�C��� ����H��� ��  P�  
 0��  S��� Y�  �2�� @�� P��  �>��� �� �@�� P��2�� �� T����,���  �  T�@��U  
(0��  S�  
( ����a �  P�    U�  
@�����  P�D�  ��� �8��	 �� ��a �  P�  
$��E � ��\  �0�����	0��0��  ����  P�%  0��  S�"  
0��	�� ������� PP�  
0��0�� �� R��  
��� R��� �	 ����$ �  � ���������0�� ����  S� ��  
 0��  S���� \�<  ��������\��������( ��,��1a � 0��`��0��e���5  �(0��  S�  
����  �P���@�� ����Oa �  P�  
 ����' �� 0��N��� PP�  '0�� ��0�� ��L��� ��  � ��} � @P�  E��� ��   �  ��(Ѝ�������� �� � `P�N��J����� �� ��P���` �v��� P�� ����� `P����
����0��  S��������4���F���F��&���F��G��#G��SG��mG�ÊG��T��+C��(C��$C�êG��EF���G��H��H��BH��{H��`��0@-��M�@��P�����  P�!   T�  ʄ �� �  � ���� ��0������  P�  `0�� ���� ��������0��0�� �� R�<�  
8 �� R�4�� �	 ��, ��0�� �  ��   � ��Ѝ�0���H��4��+C��(C��$C�úH���N-�R��0�M� ��\���  P� @�(@��  @��( �����Q �e �1p��  �0�� ���` �0�� `�� S�  ��� �� ��� ��Pc�p������� ���a �: �� �� ��0��@�����`�� ��`  �0������� ��`��0����� ���` � P� p��i  � ���� ��Pg�ia ����0z� 0�3@��  \� 0�  S�    Z�  
 ����0�� �� R�  
�����
 ��|���
 ��` ���� p�� [�J  �@0��  ��0��
�� ��Pk�Ha �@��0��  S�   ��` ���� ��� [�9  �p��(0��0��
@��Pk�@��  ���� ��4a �)0��
0��0��  S�  
 U�(  �0��r ��PE� ��o �� ��@��  ��0�� ��  �� S�  �  U�  
PE�,0��0�� `�����0�� V���  ��	p��|0�� R�  
  U�
  
PE�;0��0�� p��X0�� W�s�� 0�� 0��@��  �<0��@��  ��( ��,0�� $�, ��(��  Q� �  Q�(�� � ��0Ѝ�����4��H���F�� R��@-�`��d�M� P��@��   �����` � pP�
  ����� ������ ������ �����  � �����	` � pP�  �������� �{���" ����  P�  V�4� @�Y  "  �0�� �� R�x�  
t�� R�p�� �����p��	 �� `��\�� ���0�� �P�� �P��  �0�� 0��0��0�� ��0�� � P�� U�����`����� @���3�� T���� ��[���  P�  
���| ��C�� ��  P�  
��i��� �P�  
0��0�� �� R��  
��� R��� � ��	 ��3��  �����0�������������_ �  �|��\ �x��Z �t��t��W �p��A �`��? �d��= �  ���  �0F� S�m  �L�� �� ��_ � P�   ��T ��_0��T���  P�  �2��T��_ �� P��  �0�� S�  	0�� S�  
 P���2�� U����  � ��_ � p�� ��_ � `�� ��_ �`��`��0��  S�v`��v`��    �����  � ��_ � P�`�v`�? V���  ���� ��P��0��  \���� ��dB��d�� ��������;d � �� ��X �����  P�s  X0��  S�p  
 ��P��	�� ������ @P�  �a��Xp�� �������� PP� ��@�p�P�����  U�M  � ��������  P�   ����k���  P�G  
X �����O  � V�J   ����*_ �  P�E  @��X��_ ��T0�� ��(���  P��t�9  X@��TP��p�� W�   �����  P�*  
 ��4  ��0�� �� T�  �� �����  P�  
 P�  ��`��
 �  ��0��  �0�� �� R�`��  ��0��`�� �� B� ��   � `�� ��v��� ��D �0��  V�0C�0��  
����   �������  P�  
� ��
 �  �
 �  � ��<	 �   � ��dЍ������H���F���F��&���H��4��+C��(C��$C���H��I��,I��HI��_I�ÒI�ùI���I���I���I�Ëd���I��T���I��J��a2��5J��pJ�çJ��tJ��AJ�� R�p@-� @��P��  ��p��� ��^ �L0��  P�  ��   ��p@��	 � ��Zt �  P�  ���  ��W
 � ��p����� ��R
 �  ��p������P��0P���F-� `��$�M���P��@��p��� �  P�  
 �� ��` �x2��  �� T�  
 T�  
 T�  "  ��� �� ��` �@����� ��� ��^ �  ��  Y�(2� ��  
 �� ����  � �� �� ���_ ��1���� ��  ������p �  �O �� � ��� � @��m  �P �� � ��t � @P�P �@��d  �Q �� �1��  ��  P�  
`�����p ������ �1��  ��  P�  
`�����p ���l��� �h�� 0��  S�  
\��� �X�� 0��  S�  
L��� �H1��  ��  P�  
`�����p ���,�� �(1��  ��  P�  
`�����p ����� �1��  ��  P�  
`�����p ���� �� ���� 0��  S�  
� �� �  T�Q �  
�`����  ��]��� ��N �  P�  
���
^ � @P�   0�� �� �� ��	 �R ��9 ��� �� ��0����� @P�R �   �T ��/ � ��$Ѝ����� @�������	��H ��4�����BP�����LP�Ü3��6�ü3��TP�ü���	��p3��'��x3��]P��|3��cP�����jP��nP�� �� ��:��� �� ��7��� ��  ��4���0��  ���/��� R��A-�@��P�� `��  � ��	 ��4��p��7 � �P�  
 ���� D�0���������� ���A�� ���@-� ��c	 �  �����Q���F-� p��`�� ���M����0�����
P��  �c R�  
  �b R�"    �d R�  
t R�  
  �p��  �  S�  
c  �  S�a  0�� P�����  �  S�[  0��
P��  �0�� P�� ��  R�����J�  Z�  ����  ��- R����
P  �� �L  �@��*	 �  �� �� ���^ � Z� `� @�� 0�   �� �� ���^ � `��  � �� R�   ��  R�  
`��0��V����� ����	 �`��� ���� ��		 �  Y�  
��`F�@�� �� ��^ �  ���� ��W �0�� P�  
� ��� �  � ���� ��0'�[ �  P�  ` ��3 �\���\ �� ��X �� ���� �  � ��  �� �� ��  �8 ��� � ��Ѝ�����  S�������Q���Q��R��/R��t��p���QR�ÎR�ÛR�� R�p@-� @��   ��$��] � PP�  
 ��p@��r � �� � ��p����R���R���@-� @��P��  �= S�P��  
 �� p�� �`�� 0��@��  W����
  S�   ��
 �= P�   
 `�� �������F-� P��@��p�� ���  �	V�`��   � ��� � �P����	�� ������ �P�
P��  ����  �� �  P� ��  
P�� U�	 ��0�����:  U���, ��  � C� �  �	 ��� �  P�	`���� P�� �������R��@-�0�� �� ��t �L �  P� ����t��
S��0��@-� �
  
 ��0��  �� ���� ��Z �  P� �    �T��  �����  P�T ��   �  �����@-�  P�  �� ��  
0�� �� ��Z � 0P�@�  
 ��@ �� ��G � @��	  �  ����
 ���X � @P�  
 ��) � ���	 � ��Ѝ����'S�� R��@-�P��`� @�p�    ������ P�@�  
�/�@ �� @��' �  � ������  P�  ��@�� �� �`�� W�p������ ������.S��OS���F-�P���M����=��@�� �� `��|\ �  P��$��   3����  ��P�� �� ��� ����� ���5Z ���� p�� ��L\ �  P�  
 �����G\ �  P� �  
 �����A\ �  P�   �� Z��Ѹ�զ  ��� �  P�  � ��� �  P�  �  W�!  
��� ��-\ � P�   ��
 ��] �P� p��
  
KP�  
�P�  
�P�  
L2�� P� �D��  ��<��� �P�y] �p��z �P�u] �V � P���� Z�  �0��  S� ��p�   ��GY �Pp� P�3k  ���p��(\ �
 W� ��	�������	 ���	 � pP�	���a  
�� �����0�� �� �����  P� ����0���� �� ��
 R� ������ \�  �0�� �� �� ���Y � ��� ��+	 �  Z�  <1����8��  �� �9  � ��(���[ �  P�  @�� P�� p�� ��  T� ����
 ��   
B] �  T��  �p��T��  
@�� 0��  S�@� W����<����%<���(�4�� P��"4��0��  � ����[ � PP�   ���� ��%] �0��  ��  � ��x��[ � PP� P�  �� ��` ���m �   �P�� ��Ѝ�����A �����kS�Ä�âS�èS�ïS�öS���S�� � T���.���S��t���S���	���	��H ���	��4�� R�   �� � ���� �����@-�<0��  Q� ��  �� 0�� ��  
 0��  S��    ���� �� ���Ѝ� ���&���F-� P��4�M�p��`�� ��
@�����  �c R�  
t R�	  
b R�    S�	  
V  �  S�T  @��P��  �  S�O  
@��   �@�����0�� n����
 ��  R����`F�  V�  ���� 0��- S�C  	�����	0������ �;  � �� �� ��\ � �� `��, �� ���[ �  T�  
 �� ��,��W �  P�@���2 �  �  �,@��  U�  ��(���/�0�(@�(0�{W � `P�  ��?�� ����� �� �� �� ��� �  �  U�  
  �����/�>U �  ��@�� ��`�� ���_ ���T �����  ��  �H �� � ��4Ѝ����� �� �� ��s\ � V� `�, ���������t�À���:T�ÎR��wT���ÛR�� R�0@-�@��A�M�  �= �  � �����  P�  �  
 ��$��_ ��� ��� � ����P��X���Aߍ�0���X[��{T��  ���/��, � ���8 � ����#���/��@-� @��� ��� � `�� ��8 � P� P��� �#    �������0�� P�� �   ��? �  P�  � ��H �'  �  V�  
 ��$ �  P� ����
0�� S� �  @ ������ PP� �  
D@��`�p��@��  V����  �P������ ��n � @P�P�	  
 ����s[ �`�� ����N � P�� ��� � ���������X��V'uX�ÇX�×X�åX�õX�� R�@-�0@��  � �� �� ���[ � @���� �� � �� ��@�����  ���X�� ���/�  ���/� R��N-� ������ ��`B���@��[Z � P��p�����  P�@�`F ����  �����PZ �  P��  
  �����KZ �  P��  
  �����FZ �  P�  
  ����AZ �  P���   ���	 V�  ��  �  ����7Z �  P��  P���  � Y�    ��h��.Z �  P�   ��SZ ��p� ��3  �  ��D��$Z �  P�   ��IZ � �P���  U�  ��� �����  � U�    W� ���
�  � ��������Z �  P�    ����	Z ��p� ��3�  � �����Z �  P�    �����Y � �P���  �  �����Y �  P�    �����Y �  P� ������s  �  ��t���Y �  P�    �����Y 렯��i  �  ��P���Y � �P�  	��
 ��  ��[ �	��
 �� ��� ��[ �  Z� ����W  �  �����Y � �P�  	��
 ��  ��y[ �	��
 �� ��� ��t[ � �Z���F  �  �����Y � �P�  	��
 ��  ��h[ �	��
 �� ��� ��c[ �  Z� ������4  �  ����Y �  P�   ��
 ��  ��V[ � ��
 �� ��� ��Q[ �  Z� ������"  �  ��D��Y � �P�  	��
 ��  ��D[ �	��
 �� ��� ��?[ �  Z� ������  �  �� ��Y � �P�  	��
 ��  ��2[ �	��
 �� ��� ��-[ �  Z� ������  U�  ������ P�� ����  � U�    W� ���
��� P��`i�  V�  �	A��������  [�  
�z� ��3 z�  �3����  ����\Y � PP���
p���������i"��vY��yY��|Y��Y��6.��5.��9.��$.��*.��1.�� .��B.��&.��;.�� P�t ��/
  � P�h ��/d �5�/1 P�\ ��/ P�  
  �	 P�H ��/D �5�/1
 P�< ��/� P�    �, ���/�( ���/�$ ���/�Z���Y���Y���Y��+Z��Z��/Z��Z��8Z��a2��@-���0�� @�� �� �| ��� �� �0��0� S�d �  
 S�\ �  
 S�T �T �� ���0��H ���� �0��0� S�  ��, �� �( ��@�� �HZ��LZ��OZ��7[��zZ��fZ��nZ�ÄZ�ÒZ�Ëd�� P�p@-�@��P��  
 P�  
  P� �  
9  �� �� �  T�  
 T�1    �� ��p@�� �� �� � U�� ����
���: U�%  � ������ ��@D�| � T��  �(��0��8��@��H��P�Ð ��
  � ��  � ��  � ��  � ��  �| ��   �x ��e �t ��c � U�l ����
h �5���:P U�` ����
H ������`��� ��L ��p@��T ��Y�áZ�ýZ���Z���Z���Z���Z���Z���Z��[��[��[��"[���Z���Z��/[��<[��M[��X[���F-� @�� ��P��X � `����p�� ������6 ��� ��0��  �(�� ��  P�`� S�0������$%��  R���� 0�    �R������� \��     ����  \� ��  0���C�  \�����0��  S�����8�� �  Z�0�  � C  � ��	 � ���� �0��  V����  ��	 ��|`� `�`�� 0��
0��
���!�����0�� S�� � ��  
� �� S�� ��  �1��`��� ��0��� � ��cX �  P�  ( ��_X �  P�  H ��[X �  P�  
 �� ����(0��H��� ���� �p ����� �5��  S� `��  �  �(��p��  P�  
���� 0�� 0��5���� V�`����������W[��[[�û���_[��c[��t[��l[��}[�Í[�Ú���0@-�$�M� P�� ��  �� ��X � ����@��l���$Ѝ�0���7@-�1�� @�� S�<  !��P�����1 �0������� ���#4��  ��� �� � ��X �  P�  ( ��X �  P�  H ��X �  P�  
�� ��( ��H0�� �1��  S�  
x �� �����!������d �� �  �!����� ��P ��y ���!��D ��u �
1 � ��0��4 �����B?����,4����� ���j �>���[�ù[���[�Ëd���[���[��\��  Q�@-��M�  
<�� ��7 �@��  P�  ��� ��U �܍����H\��p@-� @��P��` ����L ��� ��P ��H �L ��F � ���� �����8 ��@ �0��  S�p��( ��; � �������� ��p@��5 �U\��i\�Õ\�Ëd�ã\��7@-� @��P��x ����* �0��l ��l ��@ ������  �  �X �����T0�� ��� 0�L �� �0��  S�  
< �� � �������, ��Ѝ�0@�� �Ѝ�0���\���\���\���\��a2���\�å\�Ëd���A-� @������ ��p������ P��  �| ����E � `��G�����  �  ��J��$���%1��| �� � V� �� �`������P��|p��1�� U����� ���A��� �d�� R��A-�@��P�� `��[  � �� ����4W �  P�  
 �� ��t��.W �  P�  _ �d��� �� �L  � �� ��P��#W � pP�  D��� �R �C  �81�� 0��  S�  ,��p�� �;  � �� ����W � pP�  �� � �� �����/  � �� �����W � 0P�%   T�  @�� ��@�� � PP�   
���� �����  T����  � ���� ��@��dX � P�� �� �� � ��@�� � `P�  
 0�� S�  
  T����	  �` ��p�� �  � ���A��* � p�� ������ ������ ��p�������g�����	]��]�� ]��\���0]��a]��f]��u]��y]�Ï]�� ��@-����� ��u Q�� ��� � �� � �� R�  
 R�    �0��!��  ��  � �� �� ��!X �0��  ��  ��� ��J � �����t0��  ��  ��9 �&4 �d ��A �`@��`0�� ��0�  S�  
&9 � 0��0��40�� 0��  S�   �  P����
� �4 �  ������������À����7��|���3^��  H8�@-��� ��! �  �����\����7���N-�P��|2�� �M� ���t��p�� ��� � W� ��  � �� �� ���W � W� ���  
 �� �� ���W � W� �� @��  
 �� �� ���W � ���
 ��� � P� `��B  ��
 ������ � 0�����(���#<��4��"4���!�� S���  
 ��� �  P�  ���� �a  �0�� S� ���	  P�� W� 0��0��  U� 0�  S�  
 ��|��� �P  �0��  S�  
h��� �
 �� �  P�X����
T��� �
 �� �  T�  :@�� �)  �`��
 ���� ��0�� � W�  �$  ��� �  �  U�  
 U�    ���� �� �	 ���� ���V �  ���� �� �	 ��0���� ��AQ �  P�  
� ��`�� �  ��� �� �`��  � ��| �@�� ���� `�� ��Z ���| ��_���p�� �� ��Z ���d ��X��� �� Ѝ����� @�����|���H �Ú���^��V'���������_�����	����O_��__�À_�Ø_�ö_��.���_���_����8@-�@�� P���U � P�
  �P��0U�. S�  0U�b0C�s0�� S� �� @��A�� ��8������@-� @�� �� ��8 ��L �4 �� ��I � ��  P�    ��0 �  �. �
 ��� � �����c`��m`��x`���F-� �P�@��`��  
.��U �  P� pj  
 ��U � p�����P��F)� `��
  � ��U �  P�    ��`��U �P��  W�  
@��	 T� ��
 ����� V�@�   
 @�� �������� ��0�� a��!��� ������|�ì�ë����N-�����M� ���`����� Y�P� @�p�K  !�� �� �� 0�� ���M�P��  �������0�� S�����pF�  �  �����0��  �� ��:U �  P����  ��0�� �� 0�� Y�@������  Z�   @�����  �pG�  W����� ���@��
�������0��p��n ���0��  P� ��@�	    W�  
 ��  ���  �@�� Z�������� @�� ��  � �����  P�  
g��� @��  ���@��( ��  �p��P��	 W�
�� ������ ���K�����`�ã`��8@-� @Q� P��  
 P�  � ��  P�  
0�/�  P�8���`0��  U�A��  
 U�8��  �P��( ��P0��,������ ��8���P���$��P �� @��P0��@���� �� ��8���  ��8���D8���!�� P�@-�  �����0�� 1����,�����D8�� P�@-�  �����0�� 1����(�����D8�� P�@-� 0����� �� ��1���� �����D8�� P�@-� 0����� �� ��1����$�����D8��0��  ��  �� ���/����0�� ���/����0��  �� ���/���� -�Ѝ��/� ��  �� ���/�@-� @�� �� �  P��� 0��@� ����@-� @P� �  
  � T� ��  ����� P�  
 ��@�����  ����� -�p@-�c�M�>��@�� P���� �� ��1���W ��� `�� ����� ��cߍ�p@��Ѝ��/�0�� �� �  
 ����� �0@-�a�M� �� �� ��@��W � P�� ������ ��aߍ�0��� -�0@-�c�M�g?��@���� �� ��1��W � P�� ������ ��cߍ�0@��Ѝ��/�@-� ������0�� ��  Q�  | ������  ���p ������l ������X0����  Q�  X ������  ���@ ������D �����(0����  Q�  0 ��@������� ��@�������`��D8�� a���7��a��%a��Ca��Ka��8@-� � @��P�� 0��  �4�����  U� �  T� ���  Q�P�  \�@�  T�  U   0��  S�4 C����  T�  
�� �������� ������  U�  
��  ������ �� @�� �� �����$0���� 0���� ��@��e��� T����  ��8���D8�Ø
�� -�0@-�c�M�g?��@���� �� ��1��+W � P�� ��t � ��cߍ�0@��Ѝ��/�0�� �� �  
 �����V �0�� �  
  ������@ �0�� �  
  ������* �@-�<@�� 0��  S�
  0��  S�  
����  P�  
���� P� � ���  ���������@-� @��p��  ��0��`�� P�)  ��� Q� �  ��� Q� �  ��� Q� �  ��
Q�  
| ��6���  � P��'U�"6�� ��:��   R�  �  ��  �L ��)��� ��0�� �����p �0����  ��( �� ���������  ������:�&�ha�Åa�æa���a���a��b���F-� `��L�M����p��@��%  � �����0����*� S�Ġ�  
 ����� S�x ����   
 B� S�  P��	0��\�� �� �� ���(X � �� ��
��� �  �8 ���������  �����
���0��pG�@��  W���� ��LЍ�����qb��Bb��]b��  P�  
0� @� �0� C�/ �� �� �� �0� C�/  ���/� �� P� �  �'���&���&���&�� ��<0��  �80�� �� ���/� �� 0��  �  Q�  0�� �����/�  ���/�`�����$0�� ��@-�@�� �� @�� ��@�� ��@��S ����8@-�H0��  P�P��@��  �  `� �� ��S �$0�� �� T�  : �� T�@�� ��8���  ��8������p@-�@��0��`��`��P`��^��P���^��P��ZE�
U�!  �  ������0��0�� P�    e����� p�   ������ �� 0b� S�  �Ĕ��� 0��  l�@��� ����
  ���`e�( ��`��0��`����Pe�P��   � 0�� ��p���`�����p@-� @P�p�� �0D� R�� ��  ���`����� Q����    P� ��  �0a� �� ������ ���� �� ��  ��0��  R�p��8�1��  ��p@�����  P����  �	  @�P��0d� ��@�� T�P� �@�P�@��@�� �    P� ��	  ���8A�� \�  0�� ��0��������  �����������  P��� ����p��R�
  *���!��@�����B��!����� �� ����)  ��� P�"��8 ��  � P�[ ��  �T P�"��n ��  �UP���w ��  �T � P�"	��| ��~ ��`���@��A���� Q�	  @��@��P�� �� �� ��  ��� Q�  
 �� ��  R����: �� ����0��0��p���`�����p��t���6���D-� ��  R�  0��  S�} 
  P�{ �@�� T�@��  �@��~T�  *����%��!��0�� S�   ��0�� S��<  
��� ������� ��0����� �����������������  
 Q�$��8��  � Q�[��  �T Q�$��n��  �UQ���w��  �T5 � Q�$��|��~�� ş���� ��  � �� ��0d� S�A�  �  S�0��  ��� �� ����� �����0��������� �� P������T�� ��p�� �� P�W  
0��0���d� \�  �0��@��0��@�� ��������0����� �� ������  \� �� ��  �0�� �� �� �� ������S�  *�1��`�����C1��p��3��0��0�����0�� �� ��-  �T�� U�#S��8P��  � U�[P��  �T U�#V��nP��  �UU�W��wP��  �T� � U�#Y��|P��~P���c��p��q����� \�	  p��EQ�����0��U��P��  ���� \�  
P��P�� S����:0��0����� �� �� ��A1��3��8�� ��  S�R  �  ���0��  
  ���0��  ����
���� �ၡ��
`�����"  �p��p��Pd� U�  � ��p��`��0�����@��P��P��`��p��@��0��0��P����������  U�P��  � �� ��0����0����P����������� \���� �� �`����
��� �P��A�4�������  
�� \����
��0����� S�  �  S�  
 ��  ���0�� ��������!��`��������
0d� S�c  �4��!�� s� p��p��p���~�p��~�p� ����� p� P��M  

 �� P�  *t1�� V�G  d1�� U�d�� ��  �� ��0�
p� p�p�3  
đ� |�T� �  b � � bP�p���>��pg�0���>��0��p�� ������ p�(  
� ��  e��0��  �� ������� V�P��p��p�� ��  
 Z�0�� �� ��  ��J������ ��
0�� Z�������� �� ��  � �����h ��0��<�� S�<0��T ��@�� S�@0��L0��0��0��0��0d� S�	  �0�����0�� ��@�� �����@��0������  ���������h��`��p��  Q��A-� @��=  � P�  � ���A��j��� P�p��@�� W�p�� ��p�� ��a��� `P�-  
��PF�<m �  Q�  
0D�  d�0����0� ��0C���� e� R�0�� e��b�P����������0��0��0��0�0� �� ���� �� �� g� R�  �0�� �� �� ��0��0�p��p����� ������  ���������
������������ ��
������@-��0�� P�� �`��p�����  U� @�� @��)  �  T�'  
 �0��D� �� Q� `�`� R� `��  V� � B�$ R�  � R�0��  � R� �� ������0��  �$ R� ������0����0� �� ��������  � ��P � ������`��  Q��N-� P�� p�� �  P�   ���N������`�� � V��E����`��`�� Y�	���@���  �$��	0����� S�  
 �� �� �� �� �  �0�   �� S� ��	���  @�� Z�  ��3�����
�f�p�����������0�0�`��`��  � Z�  � ��@��0�� ��0���  � �  @�  S�@d� �� ��M  
 S�	���=  ���0�� Z�F  �p����0�� I�$ R�0����#  � R�0��  ��� R� ��0�� �� ��P�� ��  ���$ R� ��0������P����   �� 0�� �� ��P�� ���� �� �� �� �� ��0��0��  ��� ��bP �|"��0��
�f����0�����0��0�`��`��  ���� Z�	  ��� ��0�� I�$ R���0��0����  �	��� Z�-  � �� I���$ R�0��0����"  � R�  �0�� R��� ������P����  ���$ R�0�� ���� ��P�� ��  0��  ��0��0��P��0�� �� 0���������� �� ��?  ���P �<  � ��'��� pP�Q  
0� G�0��0�� R��@���	�� .  
 I�$ R�&  � R���0��  ���� ��0�� R���0��0��������  ����$ R���� ����� ���� ��0��   �� �� ���� ��0�� �� ������������0��0��  ����O � ��b���  �
0f� �� S�  � �� ���`��0��`��0�� ��0��0��0��Q���  �
0�� ������� �� �� ��p�� ������`��0�� ���/� ��  �� �� �� ���/�x��p@-�tP��t ����� 0��	S�  �d ��p@��z���\@�� ��)��  ��O �  ��  ��D�� ��O � P���/�  ����I �0����  ��0��  ��p@��  ��Íb�÷b��, ��x��@-�D@��  �����*��� ���/�  �����H � 0��  �� P�  
@������ ����@��  �, ��@-�	�����@0��@ ��8�� S�  ����S��� S�  
 S�  
 S�  @������@�����  , ��7@-�l@����  ���/� 0��0��0!��J �  P�  �H ��:���  � P���/�  ����H �  ��  �� ��! �  �埶����� ����� ��>���, ���b�È���@-�@0��8�� S�  
S�	  
 S�  
 S�  
 S�  ����  � �����  �����   c�� ��0��  R�0�0� �  � �/�x��@-�����  �����@-� P�  
 0��! S�  ��X ������  �P ������  ��H ��M��0��L �  P�  4 ���0��0���0 �� ��, �� ������� �� �� �����*c��Xc��x��t������QR��tc��0��@-�  S�  ; ��a
 � ��@������@��t���c��  Q�@-� @��  
 �� �� ���N �  �����/�NH �0�� P�  
h �����  ��  �  �� ����0���K � @P� � �� � �
  0���0��,���, �� ��( �� ������  ����� ��Ѝ����c��t������tc�Êc���c���� �   
����0��  S�   
����0��  ���/�x���/� ���/��N-�l �� �M�@�����d!��P ��P���Pp��P`��PP��P@��P���P ��P��P���P������P������P������P������P������P������P������P��� ������� �����������p��p���`��`���P��P���@��@�� �� ����� ����� �����P���Pp��$����� ��P`��(�������PP��,���� ��P@��0�������P���4���� ��8���� ���<����P ��@��|���P��P���D���P0��l���H���L ��P ��T ��X ��\ ��` ��d ��h �� Ѝ�����;�ä;��T$��<$�� $�è!���!�ð*�Ä(���x��tZ���!�Äd��< ��X��<y���y��<s��  �� 0��0�� R�0�� 0��/�L0��  ��p@-�@�� P�� �� ��
��j �`�� ��0��F�
��i �0��@�� PP���� ��p���0 �� 0�� ��  R� 0�� �  ��/� 0��  ���/� 0��  ���/� ��0�� ��0�� �� ��0�� ���/�>���=��0�� `��/���� 0P�  
  ��@�� �� �  
 ��0��( ��  �� ����_ P����
= P�  � ��/�  ���/�H�� 0��   ��� ��0�����  R� ������/�0 ��  �������c�� R��N-�����0���� @�`�A�(    � �����S���  P�  @��  T� �����  �0�� ���q��Q��  �  ���L �  P�   ��� ��X �����>���  P�  
H ��@�����  �P��  U������ z�  $ ��@�����`��	 V����� ������0 ��'S���c��OS��8@-�<P��A��  T�
   �����0��0�� 0����@�� 0��0��@��0��  ��8���0 ���c���c��@-����  P��� ��n�������d��@-� ������  �� ��  �� �� �� ������F-� 0�� @��  S�T  
  ��  P�Q  
^  �0�� �� �� P�� S�ta�� ���lq��l�l�� � p� ��`!� 0�1�0��L �
0��0��P������ P�81�Q�����`��(Q�� V� ���   0��
 S�  1��
 S� a�  I����ML �  ���I��IL �a���0��  � 0��
 S�  
Io�� ��L � ��� ��L �	 ��� P�  � ��L � 0����P��  ��#1��2L �  �
0�����$1��%��� ��  R�h0�%!�
 �$!�L0�� 0��  ��  P���
~L �  P���
 0�� �� ��  S�  
  ��  P�  
0�� 0������  �������6�� d��<���0 ��T!���N-�p�� @�� ���+  �0����� ��  R�  
 0�����0��  [����  � 0����������0�� [�����  ��z��� 0�� 0��0��  � ��  P�  
������ ���`��P�� 0�� V����� ��i���P�� 0�� ��0��0��@��b���  T� ��	P�	`����	 ������@-� @�����  ��V��� 0��0�� 0�����p@-� PP�0�A�  p���  ���K �  P�  
@��  T������p���0��  S�H0��a��  
��< ��p@�����  ��8��� ��6���0��`�� V���� �� �� ��p@��-���0 ��,d��@-�����  P��� ���������d�� 0��p@-�  S� P��@��  
 ��  R�   0��  S�  
 0��0�� 0�� ��`�� ��������� 0��  ���0�� �� �� ���� 0�� ����  ��p���p@-� P��P�� @�� P������P��P��P�� 0�� ��0��0��p@������p@-� @��`������0�� P�� ��`�� ������ �� P�� 0�� ��0��0����� ��p����@-� `��@��q��Q��A  � ��  ��K �  P�;  0���  
 �����0�� S� S p��  _��� ������  ������ �� �� �� �� �����p��  �0��  S�  
 ��0��R3�� �  I���0�� ��0��  � �� �0�� ��  
�� �������� �� 0���� �� �� �� �� �� ����� ������ ������P�� U���  ������\������F-�0�� `��P��  S� @��  0��  S�N  
0��  S�  
��� ������ 0��  S�  0�� �	  
 �������  P�  
 �� P�  � ����� 0�� ��  �\ R� ��0�0��  S�  
  ��  R�������� pP�+  
 0��  ��  S�0������������������  P�  ��  
	q�� 0��
1�� 0��  �\ R�0� �� ��  S�  
  ��  R���� @�� �� @�����0�� S�  �� ����� ����G��� ������  ������ �������F-� @�� ���P��`��E  �
 W�P�	  
�j� ��P��������
��	 �� @�� ��J ������	 ���J �  Y� 0�� ��� 0��+  
	 ����� `P�   ��1��$ R�	   ��$b��? R�  ������L"�� `��O �  �a��  �  ��J �  P�  `��  V�  
  �`��  V�	�����
  � ���J �p�� ���������� @�� ��gJ �P��`��P��0��0��
 ����J � pP���  U�  

 ��J ��� �� �����
�� @�� ��QJ �  � 0�� 0�� ��
��J �  P����  T� �
 �����0 �ÃC���D-�!�� 0��p��0�� � p�X  
�K � P����� @P�  
l�� p�����M  � ��=��J �T1��  P� `�`�@��A��  �  ��ZJ �  P�  
@��  T������>  � ����PJ �  P�    W�2  �0��  S�p�p�.  
,  �0��  S�  
��� ������.  �  W�  �0�� S�  �0��0�� �� p����� ��oK � ��  � ��kK �  P�  ��  
 �� p��{���  �h0�� ��a��`K �p��@��@�� ��0��`��  V�������p��   �p�� ��h��� ������ ������ �P���� p������H��Bd��0 ��,d��@-�P ��G���L0��H@�� ��  P�P�� ��8 �P"�,��J �, ��������$ ��������P����@������d��0 �Éd�Íd�Òd�� ��p@-� R� @��`��
  � P��e��d0��0�� ������  P�  ��   ��/��� 0��  S� �p����  �� ��`��
 ��0��0�� ��p���  R�p@-� @��P��  
, ���I �  P�  
 ��\������  P�p�� ����p@������d���N-�0�M� @��`�� �� �� ��P��ZJ � ��`��������0� S�  
p�� �����0��0�� � ��X5��  R�0����� 

 Z� p�  
 ������ p��  Y�  
0I� S�  �(0��  S�  

�� ��@  � Y�   ����J������  P��  
 Z��   ��������  �
 Z�  (0��  S�  0��  S���! 
 Y��  
& Z�  
  �# Z�  
$ Z�0  
" Z��  �  �; Z�  
  �' Z�  �  �\ Z�  
| Z�  �  � 0��  S�  (0��  S�  
	  ����� ������
 P� p ������  � ��#��( ��{���  � w�  
p��
��( �� ��s��� ������ �� ������ ������#��p0�� ���0�� �  
 ����C��� 0�� �� �� ��  ����� ��
��9��� ��p������T#�� ��� ��z0��0��0�0�_ Z�0�  S���� ��4  �? P�  
{ P�p��
� ����  � 0��p���� �� �� �� �����
�� �����	�� ����� ������� ������T  � ������� 0�� �� �� �� ������   ����� ������ 0��} S� s �� �����} S�;   ��������9  �0��,0��  �0��  S�:  
���� ������ 0��' S� s �� ����� s�'  $  �0��,0��(0��0s� 0�3(0��  ��� �����p�� ����  � ����{���& W�   ������ ����	  � ����p���| W�   ������ �������  ����  � ������ p� ������G  �81��  �����!��#  ���� 1��  ��!��@  ������	 ��P����� ��������� ��  ��� P�� ��D��� u�
  	 ��x��� ���0�� R�P�"  � ��P��)���  � u�0�q�  �0��  S�  
 ������ ������0��  S�  | ����� 0�� �� 0���� �� ��,0��(0����� ��T��� z�  
 ���
  U� �0Ѝ�����0��  S���p��  W��������d��0 ��H��>�ád���d��@-� �� 0����0 � 0��0��0��0��0��0��0��~���Ѝ� ���>��l@���@-� @P��M�`��'  
 0��  S�$  

��LH �  P�  
0��  S�  
 ��p��OH � ��^����� P���G � ��\���G � �������� ����Z��� @�� ��g���	  �P���� ������ ����O��� @��   �@�� ��Ѝ�����d���N-� P��0�M� p��%  � �� R� 0�0� R�  � � ��  
@��  T�  ����7�����A��� �  R�  
0�� S�  0�� 0��  S�  �  S�  
0�� S�  
����87��  �����!��� �p��  W����0�� p��p��@��������p��`��p�����p��p�� �0��0C� S�
  ����#���  P���� ��  Q�P� � ����p��	 W� @�@  T�  
@��@T�@�� � W�  � � W� ��0�� �� 0�� �  P�  �   R� �� 0p� 0�3 � �  W�  � �$ �� 0��  W�{    ��  R�  
  V�Z   �� ��  ��  R� ��l 
 �����@�� 0�� 0�� ��0��G � �� �����p��(���,P�� `��5  ���� ��� ���%  �  S���"  
�G � pP�Pi�  	 ��G � p�� P���� ��������� `�� �� ����������,G ���4��:G � ��	����BG � ��1��@��P�����P�� 0��0�� 0�� ��	 ��  S���� ��0�� Z�  

 ���������� ��  P����,P�������(���0��p��`�� 0��  ��  �� ��  ��0��  R�   0�����`�����@��  ��}��� ��{���0�� �� 0��  �� � 0��  ��  P�   
q���0�� �� 0��  ��  � W��  
	 W�    [��  
  �
 W�  ��  [� �����  � �� 0��  S��  
 S��3�� 1��0���  @�� ��  P�  
����  � 0��  S� ��  �  ���� 0��
���
�����  P����  Z�1  
 0��	���  Y� ��,    �#H �=�� ���G � 0P�
 ��  �  �1��� 0��	 ������ �� ���a��� 0��
 ��	0����� Z�   
$��� 0��	���  Z�
 ������  � 0��
������ �� ���N��� 0��	 ��
1����� Y�  
0��0C�0����� 0��
���
�����  P���� �� 0��  R�;  
0�� ���0�� ���0�� @��0��(p��  ����� p���F � ���� ������  Y� @�� ��  
4��yF ��� ��vF � ���F ������
0����� W�  �� �� �� ��   
���� ��
0��  S� ����� �� 0��(p��F �
�����  �� ����� 0��0��B��� ������1��L���7  �	 ��;�� ���F � 0�� ���  P�� ��t�	   �� ������ ��� �P�   0�� ���P�������(  �0�� �� S��41�� R� ��0��� j� R�  �	 ����� ���  � 0��	 �� ���0�� 0��0������0�� ���  S�� �1� ��� 0���l� ��� z�  �� ��0��0j����L2��  �$0��  �� W�0�| ��  S�
 � 0Z�0� W�  ��L2���#  
 W���  Z�0��   S�   � S���   
���@����  Q�P�P�  U�I��
 ��0Ѝ����� �������0 ��6.�û����d��e��h���, � ���8 � ����#���/�@ ���/� �� P�  � ��/�@-����� 0��   �0��!��  R���� ����� 0��  � P��  
0��  ��  P����� ���/�  ���� ������f��\��  ���� ������f�����  ���� ������/f�ì	��  ���� ������=f��<
���/�  ���/�@-����  P� ���  ��n P� ����@-�  �����  P�  ����� �� ��@��9G �Qf��8@-�P�� @��  � ��  P�  
�E �  P�    ��8���@�� 0����  S�����  ��8���  ���� ������Ef��<
��  ���� ������h�ì	��  ���� �����������  ���� ������Wj��\��@-�  ��~���0�� P�  � ����V'@-�����  P� ���� ��q��� ��o����N-����P��`�� @��w��� ��� ��m��� U� 0�# ��� 0�% 0�%���(�� @��]���p��  ��  ���p��W��� �� �� @�� W����������@�� @������@-� @���� ����� �� �� ��@��? �[f�Ëd���@-�  ���M� @��0��P��P������D��H������ ��W��� `�� ��Z��� P�� ��]��� p�� ��`���0�� ����  ����������� ������ ��������� ��������  ��� ������ �������  ��� ������ �������  P�   �������  P�   
 �� P�����x�� `�� �����  ���� ��\��x ����� ����� ���� ���  P�  
  U�T ��,��  
 �����P�� U�0���� �� �����:Ѝ�����4���gf��}f�Îf�Ýf�îf���f���f���f���f�� P��/�E ��F-� p����P��@��`�� ������  P��� 0�  
 �� ��VF ������ 0��  T�.  
  Z�   @���� �� ��@�� @��C �
 ������  S�  
 ����*��D �  � ����*��
D �  �� 0��  S�  ` ��P���  ������ ���  �  ��H �� ��  �� ��Z���  ���� ��8�����$ ��?���  ������ @�� �� @������g��g��7g����@-�H ������ @P�  
 �� ��hF ����, ������ 0P� �  
�� ��_F � 0��0�� `����cg��Qf��8@-� @��{��� P�� ��������8��  ��  ��> � P�� ��i���  U�  � �8���0@-�D�M� @�� ��@ �� ��RE � 0���� ��@ ��0��> � P�� ��U���  U�  � �DЍ�0����F-�(p��,P�� P� ���`�� ���@����� ���  � �����ND �  P�  � �d  
m  �D0��  S�K  Z  ����������	 ��x  � ��@�����  P�  �������	 ��  � ������  P�  �������
 ��g  �P  �
 ��d  � ������  T�  
d������ �����  P�  P����� ������D����� ��R  �0�� S�  0��
 S�   �������  P�  
 ��*��� �� ����� ��@  �
  � �� ��� �� �����  �� �����  �� ��������  � ��������  P�
  
 ��+  � �� �����  ���� ��0��o���  � ��   � 0�� 0��0��0��  S�  ��� �� 0�0� 0�	 ������	�� �� ��WE � `��P��� P� ����������][��ng�����������	���æg���g���g���/�@-� @��   � �� 0��  S�	 S���
  S�  
��@��   � �� 0��  S�  S  
	 S����  �  S�  1��  � T� 0�� 0����� ����U��� �����j�� R�p@-�@��P��`��  �p@������  ��`��������  P�   ��( ��A���  �W���P��  P�  
 ��p��� V�����p���OS���N-���M� @��P������  T��  
 0��  S��  
 ��C �� P�  ���� @������  �o���� �� �� �� @��:C ��  �' Q�   S�\ P� "  R�
  �S���; Q� ��  \�  
S�\ Q�  �0�  0�� ��  Q���� ��0��}C �0�� ��������E���@��  �� ��P�� ��0��l  � Q�p��PE����R  
\ Z� ����\ P� ��  \�  
  U�a  
���PE�\ �� Q�  
 Q�  
\P��' Z�  �   P�`��p�A  $ Z� �  Q�>  
`����p��$���A  �( Z�{ Z ��`��:  
�Y�$ �� ��3  
-  �) Z�} Z��`���  �  
(  ��������� Q� �������ύ� `����DcA� ��?��� ��  P��    ��I��A�������`����  Y�  \���  �\ P� �' Z�  �  P�  
`�� ��p��'���  ��I�`�����p��  �`�� ��p��@��
 ��  Y�  U���  Y�@���KE�� 0���� 0�P����� pP�  
��e��� `P�  �� @�� ��t���  �0�� W�  ���� @��  ����0�� \�   �  
� �� @��P���  �P�� �����?�� ��<�/�`��  P� @����  P�   ��  � ��`�� 0��  S�0�  �D��0��  T�@�   � @�� ���ߍ������j��e��h��2e���D-�@�� 0�� P��`��p��  S����)  
0v�	 S�    � ��� 0��0C� 0�� 0�� ��
 S�����  � 0��  ��	 S�0��  d0��  �  ����� 0��0��0�� 0��  � 0��  �����P�� U����:  �  ����� 0��0C� 0�� 0��0C� 0�� ������
�È
��  Q��A-�`��@�� P�� ��   ���  ��  \�#   p�� B� W�  � ���A�����  Q�p�� p��  
 ��pa� W�  � �� G���  ��%C � 0����\ ��P��  �� ������ 0��0�� 0��   �j���pW� ��������� 0���� ��P��  �� ������ 0��0�� 0�������j���N-�(��� `��p�����P�� @��,���  �0��� ��@�� �����  U���
 ��	0��PE��������0���@-�0�,�M�@�� P�� 
 8��  ��  R�  �ǟ� ���� ��� �� ����� ���7�� ����P Q� 0��1������7�� ��  ��  U�  
 ����� �� 0��0��0��B � P�  
 �� ��0�����@�� ���̠�������p�� `�����p���
 \� \ P�P�	  
 ��	���P�� 0��0�� 0��! S�  SQ 
> �  V�.  
 V�  [ \���`����
�� �� ��0�����@�� ���`��̠�����������A0L� S��  �o���o���l���m�Øl�Øl�Øl�Ìm��(0������� �� ��0���N����@�� ���̠����y��������� \�  � \�Z  
  � \�>  
  � \�2  
C � \��    � \�"  
^  : \�  � \�f  
  � \�]  
 \�  
 \��  �  � \���`����
  � \��  V  � \�g  
� \��  d  ����0��0C�0��0�� ��  S��������0�� �� S���* �� `�����0��0���  �0��  S�~��
 �� `�����0��0C�  � ��P�� P�t��*PE� PU�	  
�� ����  ��/B � ������ ������  ��y���PE� ��v��� u����H  �0���� S�[��*c�����$������ ��i���0�� ��0C�0�� S�����N��� ���� R�J��*b��  �p'�F���Y���0��0C�0��0�� ��  S������  Q�;��
T��T$������ ��J���0�� ��0C�0�� S�����/���0��  S�,��
P�� C��� ��Pc� �� ���A � ��6��� ������� �����  ��/���PE� ��,��� u����0�� `��0C�0�����#��0��  S�  �C��� q���|� ����p�� ��  R�  0�� `��  �h3��!���k�  �D3�� ��  R�����0�� ��  R����
�� �� �� R�  �� ��3��#��0�� �� S�c�  
#��1���k�  V�   ��������������0��0C�0��0�� ��  S������  Q�
  
���"��Y��� ������0�� ��0C�0�� S������� ��k@ � ���@ � ��  R� ����* b� ��T��D���0�� `��0����� ���� ��0��̠���-������b���� 2�� ��1����N@ � ��0�� S� 0�� S�0��0���1�� �� �� ���1�� �� ���1�� ��k  �  P�$0�� `�  
�@ � `�� �����P�� `�����pp��
 W�  
  � W�  
 W�5  
  W����
:  � W�  
  � W�5    � W�  
 W�0  '  � 0��D�� 0������ d�D  � 0��  �� 0��@  ����� 0��0C� 0�� 0��� �� S����� 0��P��$0������  ��$0���� �� `�����$0��  ��  S�$0�� P�� �� ������ ���  \���������� ��  ��$0�� `����� P�����$0��� S�  �	 W� 0��  t ��0� ����� 0��0��0�� 0��  � ��0�� 0��F���p��$0��0��$0����� ��?������,Ѝ�����"�Ä
�ì6���j���j��a2�ÀB���j�È
��0��  ��.C�A�+C�����B���@-����� ��/���  P�@�  
 ��
 ��A � @�� ��&��� 0P�0�  T� `�� 0��  S�"  
� ������� P��  � p�����p�� PP��  
���P�� @��  �3A �d W����@D�L ����x���0u� 0�3  T� 0��  S����
 ������  U�   �������q��������j��N���j��k���F-�!����M�!�� 0��  �Q��A��� ��Q��0��  R�@��a����� P��@��  ��p��  ��@��P�  R�P�  �  
0C� P�� ��1��  ����� �� R�0C����:  ��  ����a���5� Y���� ��  
0C���1��  ����� �� R�0C����: ��  � R�p��@��0C����: ��Ѝ�����00@�s ��	 R� ���/�a0@�s0�� S�W @��/�A0@�s0�� S�7 @�  ���/�8@-� @��  ������ PP�  � ������  P���8���  ��8����N-�@��P�����  �S R� ��  
  ��0��  R���� ���  [�
`��  
p�� ������  P�  ��}  �00K�	 S��{  �lv��|v�Ìv�Üv��4x�ìv��4x�üv���v���v��0@� `�� 0��  �0@�`�� 0��  �0@�`�� 0��  �0@�`�� 0��  � 0��`�� 0��
  �0@�`�� 0��  �0@�`�� 0��  �	`��0@� 0��0�K�  ��p���p��{0��  ��	 S�J  �0��{������#2 �0� S�  � �  A�  >  � �����  P�8  � ���p��  ��z��� �����  P�0  � ��� 0��p��z�����  �� ����� 0P�&  � ���p��0�� ����� ���~���0��  P�  �������p�� ���z��� P��  �s���p��  P�p ��
���  � ��P�� 0��z��� �� U�����f���  P�  �
���p ��z���
 P�`�  �`��   � `�� ������  ���/�h��0��  ��  �� ��4��  ���/� 8�� 0��@-� @��  �����4@��  T������� 8��@-�0�� �  
$0��0��  S�  ������������������ 8��@-�0�� �  
$0��0��  S�  ������ ������� ����� 8��@-�0�� �  
$0��0��  S�  ������$�������$����� 8��@-�0�� �  
$0��0��  S�  ������(�������(����� 8��0��@-� � @��  
(0��0��  S�  ����,0�� ��3�/������,����� 8��0��@-� � @��  
(0��0��  S�  ����00�� ��3�/������0����� 8��8@-�<0�� P�� @��  �>> �  P�   0��@��8���4@��  T� ������� ��8��� 8��@-�$ ��r���  ��p��� ��n��� ��l���h���@�������
��0��h�à�À0��0@-�D�M� @��  ��> ��� ���= �0��,�� ��0 �����0��0�����$�� 0��$0��( ��00��(0��,0��3  �4@��P�� �� T�< �� �����DЍ�0��� 8��  ���/�<8��8@-� PP�@�  
 ��<����� @P�  
��< ��> ��� �� ��= � ��8���p@-� `P�<0�4@�
  
  ��= �  P�  
 @�� 0��4PD��� �� T���� P�� ��p���8��<8��@-����� 0P�  ���  ��4���  ��4��4��8��8��� ���8�����8��@-�l0��@�M�< ��@��4��� ��8���4��� ��_> �H�� ��= �1��0�� ��40��$0��00��(0��,0��00��(0��,0���������  ��@Ѝ����8��k�Øy���y��y��Xy��0�� p�  �3  ���/�P8�À ���� �� �| ��/�0�� �� �@-�0�
  @��!����� ��4��0�� ��0��4��|0����� ����.0�0� ����$��0�� R� ������@-� @�� P�� p��  �����|��0��� ��!� 1�� V�`����J������P��|p��1�� U� `������  ������H% �0�� ����� q�0�  � ��/�P8��0��  ��,)���/�(���4 ��@-�,9�� S�  ʓ������,������� ������  �����(���k��8@-�0��0��  Q�  x ������  ��8���H� �hP��� �� @��0�� �� ����� E��0�� �� ��� P�(ł� �����(@��H% �PC� ��A!�@�� �0:��(Ł�8���(���?k��P8���N-�� ��0�� @��`�� S�  
��$�����  ��������  �� �� ����= �Q�� 0��G���1�����
p��3  �0�� S�  
 S�&    ���0��
 S�  
q��|���0��1��
� ��
 �����= � 0��%1��0��&1��1��  �| ��G"�&����&��  �|0������ ��J��%1�����%��� �� � ��= �  � 0��  S�	  

0��  �����P�����E?�� ��0�� R����� ������dk��a  �,0��@-�4
��  P���  ��4*��0�� ��  ��b���@��X  �(���P8��@-� @��   �> �  T����@D�������  S�8@-� @��  ����ŀ�>  �P��  �5��  S�  �����  U� ��PE������%��0��  P�  ��8��  ��8����F-�8p�� @�Ḣ��  W� �ἒ�����  � ��  ��  R�   
����:j �P��0 �嶠��`��8:��1�㶐��`��9
�� ��5��0�����T��� ���  �  W�  
  �5��  S�  �����  W� ��pG����5��  S�U�   
 P�� ������P8��(���`���p@-�hP�� `��q@��Q�����M�P�� ��T�� ��0�� �������@�����`��� ���������Ѝ�p���0@-�h��� P���M�@������� ����� ����0�� ��������������`���������Ѝ�0���0@-� P��h@���M�q�����A��r��� ���Ą��� ��#0�� ������d��������������Ѝ�0���0@-� P��h@���M�q�����A��r��� ���Ą��� ��#0�� ������d�����������t���Ѝ�0���0@-� P��h@���M����q��A�� ���� �� 0���� ������������d������_���Ѝ�0���@-��M�r���0���� ��h��� @�������������Č���)̠� ���)�L����d������H���Ѝ�����F-��M� @��`��8���p����� P��h��� �� ��� ����������0��Č�`�������̇� ���y������d������+���P��  P�  � U����Ѝ������@-�q`��rP�������� p�� ��@�� ������� P�  � ���� ��0����� ������� P�   ��� ���� ��0�� ������� P�  � 0��  S�  0��  S� �    ���T����� �  
�� ��  Q�    R�0������ S� 0�    0��  ��  S� 0�� �� P�   �  ������H��  R�  S�D-�p���M�@�� 0�0�`�� P��0  
  Q�.  
 0�����  Q�  0�� �����  P�%  � 0�� S�"  � �� ��0�����4�� 5�� �� �� ��0��������  P�  �pG���� �� 0��	  � S�	  *�� ��  Q��?������0�� P�����  �� �� ��   �  ��܍�����0@-�hP���M��� 0��q@��Q�������P��@��T��(@�� ����0��~������@��d��� ���������Ѝ�0���0@-�hP���M��� 0��q@��Q�������P��@��T��(@�� ����0��~������@��d��� ������v���Ѝ�0���0@-� P����h0��@���M����q������
 ��!0����~��� ��� ���������d������_���Ѝ�0���0@-� P��h@���M�q�����A��r��� ���Ą��� ��!0�� ������d�����������I���Ѝ�0���p@-� `��hP���M���� ���Q��q�� ����0��	 ���� @�����������d������3��� 0P�p0�l0�  � �Ѝ�p��� 0�����0@-���@���M���  ��  �Q��|�� U�  |��2"�&!�� R�  �    � ��  R�������` ��P���  ��  �h�� �� P�� �������0��|���������� ���}��t@����� @������������� �Ѝ�0���k���� ���@-�����M���0�� ����d@�����@�� �������������Ѝ����p@-�hP���M� `����Q����P��B��T��0�� ��0����~���@�� ��� ������d����������Ѝ�p����@-�rp��0��@�� ���� P��	`�� `������ P�  ��
  �  P�  ���H ������  ���< ������  ��
  ����0��ă�\����� �� ��0���� �����������k���k���@-�h0�� ���`�����w�����M��� ����0�� P����� @�� ��KϠ�P�����P�����  P�  � V� ��w�� ��h0�l0� V�0��t`�p`�@�� �����p���p��Ѝ�����p@-� `�� @�� P��  �����	 �� ��T���5�� �� �� T�@��������p����N-� `�������� p��P�� �� ��p��������� ��?��� ���� �����  P�� ��  �����@����   �  
 �  
 ���� ������@�� ��  �(��� W����  ������s@-�P��`�� ���� @��s���  P�2  ��0�� �� ����0����� �� �  
R?��0��1��  S�  
 �"  
� ��	��� ���� �����  P�  ���d ��`���  �� ������q��� ��� � 0��  ,� �Ro�� ��`��$E�� ��1��  �  P�  
 ���� �����|����k���N-��M� @��F��� PP�|  
`�� @�� �� �������  P�t  � ���� �����  P�n  ���  �� ��L: ����0����� �� ��4��0��#4��0��: � �� �����: � �� 0�� ���!�� ����0�� �� S� �������� �� 0�������  ������� S� �� ��0������0�� ����5�����  P�=  � �����@��� p��3  �`�� ��/��������  P�*  �<�ⶠ�ᴰ�� �  
 ����h��� �  
 ���� �� ���0� S�  (5��  S�  
�� ��Y��� �  
 ���� ����� �  
 ���� ����� ����� �  
 ���� ��������p��5�� W�����  ��   �  ��ߍ�����|0��#�F/��!��	 Q�  "�� Q�  � �� R�  .��� ��  R�  �+1��0� S�   d���  ���/��@-� `���M�@��� p��0�������h0�� ��|���0����� @�� `�� ���$U��q��� P�  �0��  U�%�1��0�    �(��0�� Q�  
`�� V�����  �/��$���� ������  P�  �  ����|��� ��q  ������,  �1�� S�|0��0��
  
  � S�    �  S�  
@ S�    � 0��  �0��  �0��   �0��h0�� p�� ��&���  P���X��  �
 ��P������  �� ����<�� P��+��� P�  ��	  �  P�  � ����I�����������E�������P��  �� ����1�����  �� ��w��� ����� ������� PP�  
%��� ����0���  ��%  �`����  �� �� 9 ���  ��( ��9 ���H ��  ��9 ���  Q�  
 �� �� 0��������  Q�  
 ��( �� 0��������  Q�  
 ��H �� 0������ �� ��H���  ��ߍ�����l��@l��^l�×l���l���l��p@-�X@��\�� �� ��H% ��8 � 0��H5�� T����4@��0��0:�����F���  P�  
 ��p@������0�� ��p@������T8��(���3m��Hm���@-�\0��\@��`�� P�� `��@Z��0Z������D ������� � pP�  4 ������@j������4j�� ������ ������  ��4Z������P8��(���`m��hm�Åm���F-�   � �� ���  \����
:  �  \�
  
0 T�  ���A@L�t@�� T� ���|��x \� �`����0pL�A@L�w���t@��	 Z� ������ T� @��@��
���  apL�wp�� W�  �  �  Z�@�	  apL�wp�� W�W@L�  �  T�  
7@L� T�  ��F%� ���  �  S�  
 @��`��@��  V�  
 \����  \�  
  � P��
`����� @��  T���  R� P��  � ������  ������ �� P�0�� �� ���/���ém��@-�4 ��40��4��(��$��Ē�  P�$ ��� 4��$�� ������^������l��÷m�Æc�ým�� ������8@-�P�� @��   �9 �����  P� ��  (0�� T�@��������� 0P�  
����0��  �� ��8��蠆 @-�0���� 0��  ������  P�������l���  P�@-�@��(  
�@��4��0C� S���� 0����  ������ 0����  ������ 0����  ������ 0����  ������ 0����  ������ 0����  ����� 0����  ����� 0����  ���������0��,4�����4�/�  P����� ��@��8 �l��Ð� s@-�XB��04��  S�  
 0����  ����� 0��04�� P��`��(B����P�� 0��  �����  P�#  
0�� S�  
  � S����  � S�  
 S����  �4��0��4��k  � 4��0�� 4��g  �`��$4�� V�0��$4����� ��^  � U���� 0����  ��q��� ��V  ����x��{8 �O  � 0��l��  ��i���  P�I  
0�� �� P��$�� S�0�;�4��  � 0��@��P��  ��Y���  P�9  
0��0��A����4�� U����� 0�����  ��L���  P�,  
(4��  S�  
 0�����  ��C���  P�#  
�@��	$��4��0"�� S�  
P��� ��  �(4��  S�� �
  
 �����0 �
$��4��4�� P�
  ���0��s0��  R�P����� ������
$���0� R� �    � ��   �  ��|���@��(�� 0��  �����  P����
����l��Ð� u���v���w���t����N-� ���p����� ���@��  �4��  S�`�n  
w  �S���T2�� @P�?  ��$�� A� R�� �1  �� ��$�� �� Q�0$��  
44��  S�  "��4��$��0��S� Q�  S� Q�  0S� S�
     �4�����4��  S� ��0C�  
 P� P����
�1��$�� R�G  
4��  Q�D  
��8$�� ��8$�� R� �� b�$��;  � R�@�$   0����  �����)  � t�,  
 t�  8Q���� 0��  �����4�� S�  (�� 0��  Q�  ��C������4��0��4������ 0���� @��  ������0�� ��,$��  �(�� 0��  Q�  ��C������4��0��4��`V�P����*  T�  ��0��  �� @��$��  �xP��,4��  S�  d��
 ���� W�`��`��pf���� ������6 �$��4�� f�$��`��d��$0��  W� ����,$��  R� �  Q�d��	 ������l����D-�HA��0�� P�� �����P#�C��($��T��,T��0T�� �� �� 0��T��$��T�� T��$T��8T��4T��M���4�� S�4�@�
p�`� �0  3  ���� @P�  �0��4��  S�
  �@���� ��  R�������0��������0��04��0��  �� ��$�� ��$��  � t�  `P��pG�  W�` ��0��  ��($��07 �(�� 0��  Q�  ��C�����4��0��4��  � t�  
`V����*  �� @������l��û��à��� � @-�0�� S�  � �  P���  �����@-� @���  �  P�0�0����`0���D-� ���p�� P�� @��  �@��P�� ��`���5 ���  ��
 ��5 �  P�   ��6�/�����  T�0����� ������$���@-�0�� @�� S�%  � ����� 0��0C� S��  �\���l���t���|��Ä��Ì��Ô���d���d ��  �` ��
  �\ ��  �X ��  �T ��  �P ��  �L ��   �H �������@ ��@ ����� ��@��� �0 ��@������n�Ün�àn��*[�ån�ën�ïn�Á��ón���n�ûn���n���F-�0�� @���M�� S��i  
 �� Q��!  ꠞ��l���D���l��À��Ø��À��À���l���	��0��
 ��A���l��V��� ����������  ���V ��A0��L��  �H����V ��A0������  �4��E  �0��C  �,��Ѝ��F������ �����0��  S�  
�������� Q��  ����$���,���,���,������,������� ��   �� �����  �� ������� ������� ������ �����P��@��� �  
�t��
`�����5��uG�����u�� ��7���0Q ��� ���
 ��,Q �	��yb�0 �閠l� 0��X �� ������Ѝ�����Ѝ��F��x���?p��o��'o��Do��ao��ro�Ço�âo�õo���o���o���o���o���o�Ëd��)p���o��0����� �� ��8��<��0�����/� P� P ��/� P�  � ��/��-��M� ��� �� �� ��0����`�� P�  �1��U S�  �1�� S�  �   
  ��ߍ� ����N-�!�M� P�����@�� �� ��0��p��0���4b����`�� P�� ���  ��U Q�  2�� S�  
���"��:���o  �s?��/��0�� �� �����  �� �A   ��	 T�  � �  P�  �  R�9  
0�����0��  P�4  <�� ��0����� ��  �� ����� ��0��A� �� Q��  �ġ��ء��ġ����� ���������ġ�� ��a ��0����  � ��a ��0�����  � ��a ��0�����  � ��a ��0�����  ����a �� ��0��&9 �, �����#9 �  ��%  �  W�  
 ��  P�  
0��t���0��  P�   @�� �� [������ ��0��i���0��  P�  
 ��[���  W�0�� ���
 �`��
�� �� �x���  � �� S�0�����  ��!ލ�����Np��yp�Þp�åp�ìp�õp�þp��G��@-� �� �� ��0�� ��a�������N-��M�@�� p�������� �� ��0��`����`�� P�� ���]  ��U Q�  2�� S�  6 ��d�� ���3 �  P�N  
R ��P�� ���3 �  P�A  G  �"��8��G  ����  Z�  
  V�
 ��  
���  P�   �����  �� �� ����� 0��
 ��0��	�������	�� ������ ��0�� ���  P�� �������p���  V�  
 ��  P�  
����  P�   ���0�� T�@����� ������  P�  
 ������  V�	0�� ��� �� �����0�� U�P�����
  �u_��?��P��0��0��@�������( ��- ��F���ߍ�����Np���p���p��yp���p��a2���p���p��@-� @�� ��8��� �� ��0�� ��@��{���q���� 0�����1���� ���/�p@-� @��`�� ��P������0�� ��U��  V�0��0�0��p���  ������  R�0�� ��!��0��0�0���/�0�� ��!�  � ��/�0B��� S�0�����1��1��0���/� R�0�������1Ñ!�� ���/� R�0���/��� ����0�������/��, � ���8 � ����#���/� ��  ���/�  ���/�@-���������-�$�M� 0������� ����0�����0��0������$Ѝ� ���0��<���-�  Q�4�M��������� 0��0�� ��$0��(0��0��0�� 0��0��<�� ��  ��,0������4Ѝ� ����-�4�M�  ��0�� ����0����� 0�����0��̠�0��0��,���$0��(0������4Ѝ� ����-�$�M� ���(������ ��4�����0��0��0��0��0�����$Ѝ� ���0�� 0�� ��@-� Q� @��H0���M� ��%  �������  P�!  �0��  S�  �0��  S�  �0��  S�  �0��  S�  
0��<0���0��0� �H �0��.�  H ��0�,� �  
1.��0�� ��H �� ���� �����܍����?  ����-�����4�M�����  �������̎�80����� 0��0��0��0��$0��(0��0��0�� 0��0��@0��,0��c���4Ѝ� ���@-��������4 ��8��� Q��! Q�D�%D �5����@������@-�h0��,��� �M� ��� @��0� �� S������� �0��0���0�����0��0��?���  P�  0�� S�0� �00� Ѝ���� ��      ���/��D-����� �M� 0��p������� ����� `��>���0�����@��@��"���P�� 0P�#   ��0��>0��0��0�� ����@��0����� 0P�  u�� �� ����0��>���s����� ��	��� 0P�  
��� �� ����>���0��@�媣������������ 0�� �� Ѝ������b�燐� p@-�l��� �M� 0�� �� `�� ���� ��0�����@��@������P�� 0P�	  ������(��� �� ����0�������� 0�� �� Ѝ�p��� I� ��-�$�M� 0����� ��0��0�������0��0��0������$Ѝ� ��� H��N-����(�M� P�� ��p��P��
��@�����<��@�����<�������  W�  0��0��$3�� ���� ��$p��0��0��0����� `P�  <0��  S㊤��D�  
00���  T�  *T���!��1@�#@�3  �;��$%��#;��  S���@���@�00�� �������������� 0�#0��0�� 0�� ��$0����� `P�  00����� ��������
������!0�$0��0�� 0�� �����$0��o��� `P�   ���� ��`��$`��&0��0��0��0��c��� `P�s  <0��  S�D���  
00�����Y�����������0��d0�� 0��7��� 0��d ����� ��  �>N �  Q�  ���,���
 ����7N ����  Q�  h��$���	 Z�
 �������:<0��  S�  
00���  <�����8����� T���  � D��7 � R�  �0� �������&  �5���������� ��  � T�  �� ��������  � D��7 � R�  ����� �������0��+D� R�  ��5���������� ��%c�  �
 ��:������p ��*c�����  W�  0��0��d0�� �� ����$p��0��0��0������ `�� ��(Ѝ�����=q��Rq��eq�� I�sq�È��Ëd��{q�Ïq���q��r��r���q����  H�P0��p@-� `�� @��  � ����� 0��4 ���� S�   
���� @��P���� �� T���� ��p@�������û��.r�Ëd��@-� ��40��  � �� P�  
 0�� ��  S� ����� �����  �� ��������5r��@-�����  P� ����0��A�p@-��@��`�� P��0��i��@� Q��*  �������$���4���T���h���t��È��è ��i��   �A�� ��i��  �I�� ��i��
  �A�� ��E��i��I��j���@��  �l ��I��i��@��  �\ ��i��  �T ��A��i��E��  �D ��i��   �< ��V���0�� �`��@��p@��2 �Nr��yr�âr���r���r��s��8s��[s��Pr���F-�4�M�@��`��p����� PP� @�h  
 T�0�� ���� �� ��� ��< �� p��  R�  ��(@�� 0��0�� 0��0��<��,0��0��$0��`��@��� `P�O  
 ��@�� ��}0 �  P�F  
dp��`������� ����� �������0�� ����/ �����  �  Z�� �
@�5  
�J�1 �0�����/ ��/0�� ����0��� �� 0������  �  W� �@�$  
pG�1 �0�����/0�� �����1 � ����  �����`�� �P�  
	 V�  
���� V�  �	��` ������ ��X ��	@������(��L ������,��D ������@ ��  �< ��@������ ��4Ѝ�����s�Ês�Ös�ás�þs���s���s��t��t��+t��?t��Ot��}����F-�4�M�@��`��p����� PP�@�a  
 T� ����  ��0��0���0��<0��  S�0� p��(@�� 0��0�� 0��0��<��,0��`��`��$`����� pP�H  
 ��$�� ���/ �  P�?  
dp������������ �������0�� ��/ ��  �  W�� �1  
pG�@1 �0�����/ ��/0�� ����0�� 0��  �  Z� �
@�#  
�J�11 �0�����/0�� ���� ����  ��`����� �P�  
	 V�  
���� V�  �	��X ��h��� ��P ��	@��d���(��D ��a���,��< ��^���8 ��  �4 ��@��Y��� ��4Ѝ�����s�Ês�ás���s��bt��t��t��+t��~t�Ít�Æ���p@-� �M� @���_�� 0���� �� ��7���0��0��0�����0��V�����  ��0�� `P� ��$  0`��)���������,��� V������0�0��1�0�C��� `P����  �0 �0��  S�  �PU����*  �  U�
  �8 ��0��P0�� Q� B0 �  ��'��S/��< ��   �`�� �� Ѝ�p��� ��    @-� @�� �M����0 � 0�� �� ����0��0��0��0����� @P�  }��0 � �� Ѝ�����@-�$�M� @�������_��,��� 0�� ���� �����`�����0��`��`�� ��� pP����  �0 �0��  S�  �PU����*  �  U�  �S/��g��< ��(��P0��0 ��   �p�� ��$Ѝ�����  Q�@-�@��  ����@��  ZK � ��  � ���) � ������N-�@�� �M��� ��� ���!�� ��DP�������a�� �� �� ��  �� ���� ��������� �� ������ `P�  
��� p��@�������� P��  � �� ������$  �����������J��
0a��� �P�@ ��   ���С�� S�0��@���c� �� ����_������A��@���/ ������@��0�� �� S� ��P��p��P������ ��� �����	 �� Ѝ�����t�ü��� 0���@-��M�H0�� ��H��7��d0�� @��8�����P0��p��Lp��~��� PP�]  `��30��Lp��4��dP��PP�� ��H��h ��0��x���l0��h������p0��t���k��� pP�  
  V�`F����E  �x ��W���T �� P��| ��S���U<�� S� 1�X ��  
  : S��0�   
�0��00���0��0 �� R�`�	  .  ���� ������� PP�*  $ ��;����  
`V� ��0�� �� �����*T0���H0�<�H0� ��,����  
�� ��  ��0��`�� `����� PP�  0���� �� �� `����� ����� �P�H0�0�H0�   �P�� ��Ѝ�����       �D-�0�M�`�� 0�� ��������0�� @��,0��0��0��
��� PP� �� ��l ��/ �7�� ���� ��,P��8��0��0��1��0��0������ PP�t 00��`�� ��	��� 0�� ������,0��0��0�����������Ƞ�������� PP�` \P���� �� ���. �00��\���"  
!��  
 Q�    �0��,����S�� ��1������!�����	 @� ��:��#:��0��<��0��3  � ��<�� ��0�� (��0��<��5��;��)  �������'  �Q�� Q��  ꨻�ð��ø�������Ȼ�ø4��  �4��  �4��  �4��   �4��00��0�� ����S��� ��1����!?�������P��:�� ��D���,��#:�� ��0�� ��1��0����� 0�� �� ������Ƞ�,0�����0�����0����� PP��  00���  
 ������O  � $�� S�J  ������ `P�  ��� P��U����  �0�� ���� ����� PP��  0�� ���� ����� PP��   ������� 0P�  
� ��R��P���$  �����0�� Q�0��  �l�� P��3���  � Q�  ��0��� ������ ��8�� 4��0��<��0��  S�0�0�<0��0�� �3� P�  P�  
3��P��D0��0��  ������� �����  U�   ��y���  P� `��  H �� ��L0����0�H0��#��� PP�  0 ��H0���%  
�  
�7����� �� ��
��7���8�����0��p��,`��p��
���  P�A  
�� �� ����0��p�����,`��0������  P�5   �������H0�� � ��E  
B  ��	  
 ���� ��0��+���  P�#   ����$  ��	  
 ���� ��0�����  P�   ����  ��	  
 ���� ��0�����  P�   ����  ��  
�� �� ��0�����  P�  
 P��B  � ����k���H0��a � ��  
`��,�� �� ���, �  P� ��  ��������� ��O���0�� `�� ��`���� ��0��`��p�����t���l ��{0�����4��"$�� �� ��1 �p���l ��� ����\���,<�� ���\������������1 �t ��� ����R<��".��1 � ����� ����ʤ��   �P�� ��0Ѝ������t��    "  0  @   -1?  �t��#u��su�æu�� u����u��@x}�s��v�À��v��'v�æ���p@-� @������ PP�   ��������� ����� ��3��� PP�   ����� ������ p�   ��>���  P�P�   ��p@��1��� ��p���p@-� @�� ��?���0��  �� ��  �嚔��  P�  � ����� @�� ��v��� `P�  
���� PP�  
 ������ P������H � �� ��H ���@��  �� ����� T���� ��p�����ä
��2v��X0����T���@-�  ���� @��D�� ����� ���� ��0��0��	���$0��  �� �� 0��@�� @�� �����
��ܰ����è���p@-� `Q� @��  
0��
P�� ��0 ��  ��r ��(��  ��"��w���0��"�� ��"��  �  U�PE�  0 ��p@������- �0�����, ��2�� ����
0��0��(`��p���Hv��8@-�(P�� @��D��0�� ��0������ ������ ��@��(0�� Q�0�  
 Q� 0��0�0�(0��8����D-� @R�P��(p��  0�� ���   ���
`��  �  V�`F�  l�����T  �O- �0�����$ �� ����  T�  
 ��. ��  ��`������0��  ��( ��� �( ����0���� ����q���� ��0��  T� �� ��  
 �� S�0��'0�� � ��0��0�� ��
0�
 S�c ����0�  
 �0�   �0�0� � ��0� �0�  T� �� 0��0� �� 4��0 ��s0��0�� `���� �  
  T�0`��  
L  �Q����0��,  ��  
�� ����F���  ������0�� �%  
��  
 ��0���� �� S�  ��0�� B��� �� ����A�  � � S�P�����  � �0�  
0�����d ��$ ���  �, �Z����� �����  �0��0��  T�    �0`��
0�0�  S�0�����
	�0`��  
��< ��������� �  
, ��������, �  ������ ������jv�Õv�÷v���v���v��w��@-�p@�� ��l����(0 �d0��#��X2��\0��<3��X0��@3��T0��D3��6��\2��3 �|2��@0��d2��<0��h2�� 0��6��00���5������  P�  �������w�Ø���@���������À ���  S0�� ��p@-� @��/ ��dP�� 0��(0��  �  U�PE�  $ ����p@������w, �0�����/0�� ����p���#w��@-�(@�� ������0�� ��?��0������0�� �� ����4 ��8 ������  ������ �� 0�����/�0�� ���/�0���� 0��  ����0���/�7@-� PQ�6�� @��0��  
�� ������ �� ��, ������ ����, ������ ��,������  P�  �0��0C�0��0��  S����  � ������ ����, ������ ��d��, ������ ��,������  P�  �0��0C�0��0��  S����0��  S�  $0��  U� ��  ���Ѝ�0@��]���Ѝ�0���   �����c��Ew���@-� `Q� @��E  
 ��P�����1����Lu��1����� V�`�!�F �W�����F � q���� ���F � P�  � ���� �����  �P��U������ �� ����� �� ��, ����� ����, �����2��0�� ��,�����  P�  �0��0C�0��0��  S����0��  S�  @ �����,�� ��p���, ���� ��i��� ����s���,`������ � �/ u   �aw��D��p@-�  Q� P��(@��  
 �����@�� Q� ��  
 Q� �  
 Q� ��  
 Q� � �   ���� ��C��� ����t ��   � ��=��� ���� ��p@��8���  0��p@-� P��  ��d@�� ��  ��  �  T�@D�    ��p@������+ �0����� 0�� ����p���w��8@-�(@��l��W� ������� ��p �� �� �����  ����  U�
 ��PE��%  
j+ �H�� �������������0��dP��  �� ��  ��  �  U�PE�  X�����  �V+ �0����� 0�� ���� ��dP�����0��  �� ��  ��  �  U�PE�  �����  �B+ �0����� 0�� ����L�� ����������0��
T� \�L ��@����0 � ��2���������� �� ��D ������ ��$ �� ������0�� ���� S�<�<� 0�����0�� ��l��d �� ���ˌ� ������ �� �� ����� ���� ����� �� �� �����0��  ��  �� ��8���w�àw���w���w�� � �� �� �N-�`���M�P��(@�����  �  W�pG�  ���<����  ��* �H�� ������������ ��D�����  P�  
 ��D�����0�0 �  S�  D�� ����� ����"��� �� ��D ��v���  U�B  
 ��hs��9��� ����� ���1�� ��0��  Z�
�� ������� �� Y����B!��  �y��� ���  ��v��� �����
��	�R!�� ��� �� ���Z������p��j���0�� ��  ��$��  ��  �� �� �� �� �� �� �����  ��  � ��X����I� ���  ��T�������� ��0����� �� ���p��8�������0��  U� ��p�( ��  
� �� W�|��|�� �{�0��
 �
 R�i  
 �  
 �@p��p� � ��,��|��������  P�  ���������
��, ���� ������� �� 0��D�� p��0�� �  
  U�Dp��  
  �S����������Y  � �� R�) RU  
7 R�V  R  � �  
�� ��d�����4  �0�� �  
 �0�00�0�  
<�� ������8�� �� ������4�� �� ������0�� �� ������ ��  U�  ,  �Dp��>�0�  S� �����
�>�0�  S�Dp��  
��� ��k��� �� ������  ���� �� ����� �� �� �����  ��  � �  ��x ��X��� �� �����  ���� �� ����� �� �� ���������) �  ��   � ��Ѝ�������$ ��B�������x��Bx��@���gx�Õv�Üx���v���x���x��8@-���2�� �� ��@�� P��c- �x0�� �U��p ��8��l0��l9��h0��p9��d0��t9��6��8��"���9 �8��L0����8��D0��8�� 0��:��80��`:�����  P�  �8���y�è���@��Ø���y�������������À ���  U q�    ����\0��0�� ��  S� 0�0�� R������  � Q�	  �,0��1�� P�  P    S� � �� �   0�� ���/����Ü0��0C�0��  S��/� �� ��������'y��=y��$��<���@-�!��  R� ����0��  S�  
  �� ������ ����� ��1���������Gy��0��@-�  S� @��  D �� ��@������ 0��8��!��  R�  A�� ��$0�� �����0��  S���� �����'y��=y������p@-� `�� @��LP�� ��1��  S�
  
 ���' �  P�  ��  P�0�0��0�p��  �@��  T���� ��p�������0�� 0��0�� ���/�P���0�� 0��0�� ���/�P��À�������/�H0�� ��(�� 0����  ��  ���0��
�   R����*0��  ��0��P��P ��` ���/�P����N-�`��� ��P�� @���� ��4 ��E �<���2��0 �� p�� �
�� ��E �  ��
������ U� p��  
x9� U�  
  U�  D0��0#�D0��!��D0�� ���  S�������  
@ ��0�� ��0��������`��' U�@��&a��$A��M  
  � U�  
 U�1  
  U�  
Q  � U�  
  �q U�L  H  � U�@  
� U�G  @  � P��  ������P�� U�������=  �0�� �� P��@!��  ������P�� U������� @��  �~�����@�� T�������  ���P��{��� U�������"  �0�� �� P��@!��   �q��� U�  ����P������ @��  ���@��g��� T�������0��  ��@!��  ��� ��  ��� ��  ��� ��  ��� ��T���  ������P��Ô���Q� 0��4��D ��   0�� R� ��@0� � �/� �� R�0� �� � �/�P���l ��@-�8��  ����0��  �  ��A�  0S����*0��0 �� �P ��   �  
` ��0�0�  S�  
/��� �����  �����P����@-� `��  ��@�������P��  P� p��  �����
������ 0�� �� ��  P�������*��' � �� p������ 0�� �� ��  P������� ��' � 0��,��h ����,������X�� �� `����L�� ��h��D��l��@��T��<��X��8��\��4��P��0��`��,��d������P���  ������������ ��ô���4���,���p���H���@-������0���� �� ���' �  �����@-���z����� ���� ��w' �  �����0��p@-� @��`��00��6c��  � 0����������� 0��0��00���  
��0 ��C��� 0��,��0��P ��@�� T� ��P�� �� �����:p���wy��P���A� Q�8@-��� P��6���0��!���� 0��  � ��0 ��  �  
  � ��  ��  S�0C����0��0@�� �P@��  
` ��0�0�  S�  
d ��d�����0��I ��0��0��8��� �  �  P�8��< �� ��0������ �8�� ���� ������ ��8���4���P��Õy��t��íy���y�ô0��p@-� @�� 0��  �� �� P�� ��Pe� U�p��  � B� U�  p���| �� U�0�  �p��V �� U�p��U�
  �� T� �  
� T�   ���� ��  �� ��p����P�� ��$ ���������� ����p@��6���P���� B� �y��01��@-� 0��  �� �� @��!�� @d� T�  
  � B� T�,  
 �� T�.  

T�  !  �� �� T�  
  �� �� T�    �� �� T�  ��� �� T� �	  ���0�� ��  �0��� ��  �0��  ��  �T��@��  � ��  R�  
  T�  0��p ��  � T�  0�� ��  � T�  0�����p ���������������p@��  �� ��x���t �����P���� B� � �� (z���F-�P�� �� 0�� @��`�� ��0��, �� �  � �  
 0��'�� 0��  ����P���� ����T��0�� �`��`� � �  
�P��p��0 ���B � �� �� 0�� ������� �� 0�� �� ���0 ��6`�� F�	 �������� `�� �������	 ����� ������T�� ��Ѝ��F������P���0�� ��0�� �� ���/�0��"Ƞ�r �� �� ������/�p@-� @��P�� ��������  P�����!�� �������� ��������  P����� ����p@������p@-� @��P��`�� ��������  P����� ���� ������ ��!�������� ��������  P�����p���p@-� P��< ��`����� @P�  �p�� ��< ���% �d��`�� ����� p� ��   
1�� P� �<  P�� ����� 0�� ��  � \�  
� ��!��0�����  \����,  � ����8 �� ������� `�� ������?� p� V    � ��c���  ��p��� <�� ��0��&4��`��0�� 4�� ��0�� ��T ��0��P�� ��  ��H ��, ��D ��$ ��@ ��( ��< ���) � ���5 � ��p���( ���������!Ce�dz�È�����Êz�ð��Ü��ì��Ñz�Ùz���@-�@�� P��*��p�� ��f��� �� �� ��b���0��@�B@�Q `��DA��  � ��`��Y���  T� �� ��@D���� ����K���P��  P����
 ��H��E��� ��� �  �  P�  
P����L��L ��L0����D@�� ��< ��0� �@� �,��� @������[���  ������a2�ùz���z���z���z��{���z���F-��0�� @�� P�� p�� ��|�����P��P��  P�  U����&  � ��|�����P���  Z�  
@�� �����l��  �� ���Ph�� P����� ��	���*���  � ����J�	 ����� �� Z� �����	�  
��4 ��#���  �$0����  ��7 �
 ������ �� ������������<-��8{��e{�Ñz��p@-��� @������ �  
 ��d��  ��
P������   �% �PU��� ��  :���� �
 �����
  U� �  
 ��\��  ���_������ ��t�� ������   �% �PU��� ��  :����  P�
 ������  U�  < ��p@������ ����, ������ ����  ����� ���� ��p@�����x{�á{�� ��(P   p����p@-� @��P��`�� ������� ���� �� �������#��+�� �� ������� ������� ����p����@-� @��80��S�������� ������� ��|����/ ���  � ��+��|���\��X% � ��)�� ���������R% ����! � ������ �� ��,������PE����G% � u�  
 ����k��� ���� ����A( �z��� ����b��� ���� ����]��� ����
� ��   � ��P��x������ ��0����p��`�����8�� ��4��d��0��,��]��� �� ����Y�����h ��c��� ��t��'��6��� ����L ��2��� ��p�� ��.��� ��l��  ��*��� �����"��B���  ������{�à� �{���{��|��'  @-�80���� �����? �(0��  � �� @�!��0��r ��  ��0�� ������������( �40�� ��@-� @�� @��0�� @��0C�  ��0��E" �  ������ ����� �0��  Q��� 0�� ��/� �8@-� P��  �����  P�  
 ��8���0�� �� @��@������
0��  ��8��� �0��  ��  ��/� �  ������  �����  ������  ������ ������ ����� ������ ������ ����� ����� ������ ������ ����� ����� ������ ������p@-� @��P��  ����  P�p��,0�� ���� 0�� ����
0��
 T� @��p�� ��p@����� �  ������������������� ������p@-� `��P�� @��   ����� ����@��  P����p��������������������� ������H1�����F-�  ��T��� ��X@��P�� \� �� ��	p�� ��`�� �� ��� �� � P��.P��@��@��P��P��	@��@����@��@����
 �������� ���� � ��  ��0��\���` �����?���,������)��� ������`��������p����� ��� ���C���!������"���~���+P��&���,@��.��0���p���� ��`�� �� �� ����# ��$P��%@��'��(���* ��-��/ ��1 ������X���0��T ��  P��@ ��/�X��� ���/� ��0�� ���� ��'�� ��'���/�  [  0�� �� ��0��0��  S������/�  H0��' �� ��$� ���/�  H0��0��0� 0���/�  H0��(�� ��(���/�  H0��(�� ��(���/�  H ��0��T ��'�� (�� �� ���/�X���  H 8�  ���/�@-���������  ���������  P�   0�������/� P�)�0�"�0)��/�  H  P�   0��)��"��+���/� P��0�P��/�  Hp@-� 0��  ��  �@��`�����0��P��H��L�� ��@��D����� @�� R�����p��� Hp@-� 0��  ��  �@��`�����0��P��H��L�� ��@��D����� @�� R�����p���  H@-� 0��  ��	  �0��� ������ ��,L��@C�,D��,Ƞ�@C��C� R�0��������� 0H1��C0��0C� S��?  �,���@���d�����ì������������0�� ��G��F ��(  ��0��G��F ��$�� ��	 R� ��) ��  �0��B0�� S��%  ���Ð��Ü��ä��� ��   � ��x0��  �  ������ ������`0��B �� �. �  
 R��// ��H ���/�80��! ��G��F ��$��H �� ���/�0��( ��G��F ��H ��$�� ���/�X���d0��@ ��  R�  
 R�    �B�� Q� �  �B ��  R�  D����  
 Q� �  
 Q� �0��  ��H ���/�X��Ì0��@ �� R�
  
� R�  
� R��/� ��#��H�� �� �� ���/�  �� ��$ ��  �D �� �% �H �00��D �� � R�% �H �0��D �� � R��/% ��H ���/�X���p@-��@��lP��p0��x`��P��\ ��Pf� U�  � �������\�� �� ��!3��"9�� 9��:���x ��\0��0��x0��x0�� 9��  S�����p���  U�  
 �� ��������\0��H ����!3�� ��"9�� 9��#���x0��P��xP�� 0�� 9��  S�����p��� ��0�� )��p���X���  H  �0�� ��p@-�l@��p��4)��@��@b�  T�x ��p���\`�� ����= ��� P�� ���= � ��  Q�� �P� U�%f� �������� ��0��\ ��0�� �� 9��p���X���  H ��0��  ��#��  �� �� S�����/� H H0��  ��!#��  �� �� S�����/� H H00��  P�@ �,�@��T �` �X�` �X �T�\ ���/�X���D1�����F-�  ��T���@��XP��  �� \� �� ��	p�� ��`�� �� � �� ��P��P�� �� ��	P��0P��@�� ���
P��P���� @��@���������� ���� � ��  ��0��\���` �����?���,������)��� ������`��������p����� ��� ���~���&���+P��,@��.��0���p���� ��`�� �� �� ����! ��" ��# ��$P��%@��'��(���* ��-��/ ��1 ������X���0��8���0�� 0���/�  H0��  ��t ��d ��h ���/�X���0��  ��x ��l ��p ���/�X���0��| ��  P� ��/�X��� ��0��P �� �� ��' �� ���/�X���  H 8�@-�a���L0��L@��  ��H ��D0��8��0��8��0��8��<��$0��4��(0��<��1��Z��� 8��>�� 8�����X���  H  �D-�| �����x0�� P��h`��d@��`��
pF�  �����4��6��  S�  L �����
P��uP�� T����:	 V�
0V�$��r �� U�$ �  
�� �� ��� ���D������|��X��È��à|�ð|���|��p@-� `��0 ��P�� @������  ���@������ T� ������ ��p@�������|���|��>V�� �@-�@��  
 �� ��L ���  �D ��K���@0��  T��	��  
T�>�BA���� ��  �����0�� )��!#�� )���������  H	 P� ��@-�  �  
  Q�   ������0��  ��H �����(���4���X����1��p@-�1��  S�  �Q��, �������`�� ��  ��Q�� ������� ��4`��A��H0��$ S�_  
  � S�Q  
  � S�)  
 S�-  
  S�p��   �  S�J  
 �1�1U  :" S�I  
# S�p��H  �) S�'  
  �& S�G  
� �2H  :' S�E  
( S�p��  �. S�,  
  �, S�p��  �/ S�(  
� S�p��-  �F����p@������� Q� �� ����  ��� Q� �� ��  �  � ��p@������� Q� ��  � ��  ��� Q� ��  � ��	��p���p0��  ��H ��p���$ ��   �+ ����  �X ����  ���  � ��	  �G��  � ��  � ��  � ��   � ����U��� 0��H0��p���X���T��Ø�������@-�$1��@ ��  R�  
 R�    �B�� Q��  �B��  Q�
  D������  
 Q��  
 Q�����0��B�� Q�)  D��  Q�&    R�$  � ��E0����0C�p��P���� S��  ����� ������(���h0��(��p �� ��  �T0��(��p ��  ��  �@0��(��p ��0 ��  �0 ��5����� 0��(��p ��@ ��(��0��  ��H �����X���  H��� �@-�@��  
T ��@������M���H0��  T��4	��  
?��T�0���A����� �� �����0�� )��!#�� )������|��  H�0��@-�)��(!��$�� R�  &!��%A��$���'��(��"��$��!A�� ��,�� ��� ��#����  R� ��p ����l ��x ��  
R�'�# #��0�� ������0��  ��h �����X���\ ��\0��@-�0)�� ��x��(��l@��p���(��  b� �� ��x ��  R� �$#���R�'�# #��0�� ��@�����  HX��� �@-�@��  
T ��@��~������H0��  T��T��  
?��T�0���A����� �� ��g���0��@+��!#��@+������|��  Hh0��@-�d@��P;��t���8��d��h ��8��a�c� ��t �� 0�� R�  ���@������4���h ��0��d��
 B� ��$3��@��L���  HX���7}��p@-�@��~/��J��&���%Q��(3��$��Ƞ�'���Č� ��� ��d0��̌�t0��h���U �t ��d0��~��h ��0c�t �� 0�� R�  ���p@�����
���h ��0��d��
 B� ��$3��p@��"���X���7}��00��h ��,0��  R�P;��  �8���! �8�� S�   L����������X���  H|!���A-�H0��  S�Y  �p����0��`��@����� ��P��@p��C`��GP��D@��E���F ��A��B0�� Q��F  � �������0�������0���H�������0��ü���l���������$���� ��  ��T��H ��'��2��� �� 8��0  �� ��3^����������`@��\���0��2��AŌ�@��"Ɍ�|@��"9�� @��H@�� Ɏ�@;��I���  ���p@�� ��  �����3�������� 0��H0��  ����  �H���  ����  �`���	  �" ��  �  �� ��1��H��  �  ��0��H ���A������X���  HX0��X ��@-�P������a�Q�<0�5  �30�0 !�543��  S�  
 0��  S�  
��3�/� ����@�����  HX���x���@-�, �� ���(@���� �� 0��  ��;����� ;��!3�� ;���������  H�0��@-�(�� �  
I�� �   
����0��I������	  
K�� �   
_��� �   
����0��K����� �  
()��()��0��  ��� ���\0��!��  R�8���@��������H+��H+��0��  ��� ���0��1��  S�  
@�����@��(���  HX���@��� ��<0��T��)��  Q�+��()��H+��  #�� )������#�� )��!�� +���/�X���  H@-�d0����� ��  P�  
 P�  h�������D0��1��  S�  
  �4 ��"���  �����l���   �j�������0��8 ������ �����  HX���w}����Ä0��@-�@��
�@��  �  
*�� ������  ��
�  
P0��*�� ������  P���  ��  T�00��!��  �� ���0�+�  � ����o���  �����  H����@-�@@��0�� 0��� ��� ��(0��0�  S� ������� 0��0��  P� ����  H 8�@-�@��2 �� �,0�� 0��7�  
  ��@������ T���� ��@����������  H�}�û}��p@-�80��8@�� P��
 ��R��?� 0��0��0��0��0��m �
 ��P��p@��i �    [7@-�t0��t@�� P��'��<�� ��|P��'��T��HP��LP������Z�������a��� ��f���0��Q�� S�  g���
 ��N �j���o���  � �����  ��>���  X����}��@-�����0�� ��  ��!�����X���8@-�L@��83�� S�
  @S��  U�8�� ��� � �� ����� 0��83��8���  S�0�@+�#�@+�8���X���  HH0��@ Q�@��@-�@��D�� ��@��8#������  T�    �r���0��83��  S���� �����X����@-�P�� @������0�� ��L3��0��P3����� pP�0�T3�  
6n�� ��  �� ��> � �� ��� P�  �� �� ��c �Tc��L0����X �� ������PÓ�.��\#��X#�� �����TÓ������4C��������" �  ������X���~��~��~��~��$~��00��  ����0��@ �����  \� �  
 R���� 0�� ���/� ���  ���/�  ���/�  ���/�  ���/�  ���/�  ���/�  ���/�40�� ��  R��/0��!����  ��  Q� �0�� � S�����/� ��Ø����@-�@�� S�  ڈ ���@������@��p�� `�� R����s0��P��`��@��@��@��p��`��0��$��� Q�  �� B�� ���� �P��!������0�� �� ������ ���5~���N-�@���4��p���M�`��� �� ��  R����  !_����0�0�� U����� &�#�00�㌔�� ���������0�� �  0�� �  
h�����c  �0��  S�  9�� ��0��  ��}���u0�� ����������0��  �� 3��0�� 3��  U���  
 U� ��	��  
 ��� �ʠˠV=���� S� ��  ��:� 0����0��7�����V4����� U�  ��3��	���0�������� ������	  
 U� ��  �>���T�0����AI������  �  T���  
�>���T�0����AI������. Y�  �	��0 ��0��[���#  �#�� �����0��`�帐������� ��@��  �  ��)���  ��  P� ��@��  �2�帰��>������  ����	 [� ������0��@��  S�  
�  
1�����6���  ��  � S�>  
0��0��0�� S�  
 S�7    �X"�����0��  S����0� ��<2��� ��  R� ��  � ��  R�	  � ��  R�  � ��  R�!��� �!� ��1������  ��!�����0��  S����0�(���1��� ��  R� ��  � ��  R�	  � ��  R�  � ��  R�!���  �!� ��1��������`� ���h0�l0�0����1�� � � ��"���� � �  T�41��  �� p� U� ��%  
 U�C  ,1�� P�� V�$�����  �  U�z��JD�P��
 �  �	 ������*�� T���0������  U�� ������ �� ��  V�`� `� ������0��� ��  P��0� �  
  � 0��8����� �����  T�0��  ڈ���  V�0�� �� ���� �����0��l���  �� V�d ���� �����$0��� ��  P�  �0�� �� ��   �  ��Ѝ����� ���L~��l~�ï~�Î~���~��  �  �  �  �  �  �  � ��90�0 � ���/�mN�AP�  �3�/1	P��3�/1P�
�3�/1P�
�3�/1P�	�3	�#�/�`����N-�  \�5�M� ���@��l ��	  
 �� �� ��A?��<�/� P�  
��|��]���  ��(	 �3��U S�  3�� S�  
X��O  �	 �����/������  P�  <���� ��I�����#��3��$��D���#��
���4��?7��")��  S�\ �� �\ �h���  P�p ����2  

��b���  P� ����,  

��\���  P� ����&  

��V���  P�d ���   

��P���  P�` ���  
��J���  P� ���  
��D��� @P�|�  

��?��� �P�l�
  

��:��� PP�\�  

��5���  P� ��  D��������<�� p������	��� ���\ ��$������ ��*��p ��� �3��  W�p ����p`��%����#���k� � ��)����=�� ��0��  
9A����0C��/� S���� �剒��\���R㩐�� I�i6 �0��	S� �� ��  �� ��  � 4��( ��)0�� 8��*0�� <��+0��  �)<��(���+0��)4��)���)0��*������ ��d�� �N6 �l��� �����  ^��� ��0��4��  W� ��!��%�� <�� ��0�� �� 0�� ��0��
 ��3 ��0��0 ��  ��0��0��	���0��0��0��0��0��0�� 0��"0��#0��$0��&0��'0��,0��-0��.0��/0��10��20��6 ��3 ��30��8 �� ��40��9 ��_ ��L���E �� ��50��F �� ��70��T ��:���;0��<���=0��>0��?0��@0��A0��B0��C0��D0��G0��H0��I0��J0��K0��M0��N0��O0��P0��Q0��R0��S0��` �� ��U0��V0��X��\���d ��g0��W0��Y0��Z0��[0��]0��^0��_0��a0��b0��c0��e0��f0��#   ��o������� ��� ��k������� ��� �ᄐ��f������� ��� ��b������ ��� �ሐ��]������ ��� ��Y������ ��� �ጐ��T������ ��� ��P������ ��ᐐ��l �� 0���0����  P�q������0�� ��R$��� ��h�����\�������i �����.������j��� ��p ��� ��k�����Q�����l �� ��R(��� ��m�����,̠�����n �����~�������o��� ��P��� ��p�����Q�����q �� ��",��� ��r�����|�������s �����^������t��� ��P�� ��u�����!����v �� ��"&�� ��w������0���0��,*��� ���������  
 ���0��� �� ���0��� ���0����  ����<����� 0�� 0��I������ 0������ �����< �� ���4���n�(������< ��(���0��0��80��t0��0��0��x0��@0��0��h0��0��,0��$0��D0�圐��� ��  �� 0��0��͒��'��� ��� ��  ��Ȓ��"���� ��  ��Ē����� ��� ��  �㿒������ ��  �㻒����� ��� ��  �㶒������ ��  �㲒����� ��� ��  �㭒������ ��  �㩒����� ��� ��  �㤒������� ��  �㠒������ ��� ��  �㛒������� ��  �㗒������ ��� ��  �㒒������� ��  �㎒������ 0�� ��� ��1 ��!��	1����
1��*��1�� ��� �� ��W ����< �� ���0B�P��0n�DP��P0��D������T`��X���|@��Hp�����  �\ �����( ��`��@@�P�� U��  U�@��p� � 0�  0��4��	S�0��p��������`�� �� N����+ @� ��0n�@`��@��0�� �� ��l��  Q�"  
  U�   �� �� 0����� �� 0�� �� 0��  P��π���� ���Lŀ���
\��������������� �� T� 0��@d0@l 8@�5 @�3  �8���  ^�@n�  ��8 ��	 U�  � �  
�����0����  �E� Q�  � U� U    �)E� Q�  �1 U�  �����0��n� ��@��$��`��p�����0�� ���� ��$�� p��'����� U���'��`���F��'��@����*����*����*����&��	��&��
��&����$����H ����  U�  t��  S�`�������t��xp��h@��  U� ��"4��0�� 0�0�0�����P�P��0� ���,0�����4 ��0�����,0��	�����4 ��\�� U�V���l �����  R�T`��X���|@����Hp��P��D����  
0��	S� ���  ��@������@������������� ��������0�� ��X0��0��T �� ��D0��	0��P ��
 ��H0��0��( �� ��80��y0��4 ��A����B����L����N����X ��@��#��T ��@��'��D ��@��+��P ��@��| ��H ��@�� ��( ��@��� ��8 ��@��� ��4 ��@��� ��1��A��A������B��B(����!��L$��LȠ�!�����N$��N��!�����X��A$��!!��A(��"!��T���L$��%!��L(��&!��D���N$��)!��N(��*!��P ��H ��H���@��@Ƞ�B$��( ��P ��N��( ��H���@��8���D ��B(��8 ��( ��N��4 ��T���@��4���8 ��B$��X ��I$��N��4���!��I(��-��	 ��!��I,��.���
��!�� ��!�� ��!�� ��!�� ��!�� �� !�� ��$!�� ��(!�� ��,!�����| ��0��/!�� ��P��� ��1���H���2������4��3���D��5��(���6������8���7��T���9���8���:������<!��;��X ��=!��4���>�������?��� 0��e��� 0��P��  

P�$�L �  

P�ĠL��  
	P��L��  
	P�L���L��L ��P�L!��L���,$��M!��,(��N!��,,��O!��	  
+��0�� ��@1��B<��C1��B4��B(��A1��B!�����, ��0��0����� �� ,�� 0�� ��#,�� ��#$��#8�� ��0�� 4��0�� 8��0��.4��0��.8��0��.<��0��3��� ��9��0�������t��  Q�  
 �� ����p0����d�� P�a 
�� �����] � �������  W�  � ����*��`��{ �,���$���
������@��  ��~����(��V�Ä�ß�û�����������2���N���n��Ï��ñ���ƀ��ހ��������e���=��Ä��è���Ł�È��Ëd����������� ��  \� �� ��N  
)�� \�v0�� 0��B����B��B(���� ��C  
)�� \�0��B����B��B(���� ��9  

)�� \�0��B����B��B(��	��
 ��/  
)�� \�0��B����B��B(���� ��%  
)�� \�0��B����B��B(���� ��  
2)�� \�0��B����B��B(���� ��  
6)�� \�0��B����B��B(���� ��  
b)��0��B<��0��B4��B(��0�� ����� �� ��0������d����� P�  
�� �� ������`�����0�� V����
@��	���,���\ ��0@� W�,  
 ��*��d ��� �h��d0��)a� ��  R�`�����`��~!� BB�b��-�A�-�A �B  �  �    ����� ��  R�����!�� �� ��!�� ��!�� ��  �  �� ��  �� �� �����0�� \�����R  ����*��d �� �<0��h���  ��h��� `�� l�  R�0��0��~�AB ���2��$0��0�,0��d0���A��A�B�"�� �� ����� V�  ,����������  \���� Ġ�  ����� Ƞ���� ̠����  � ������ ������������`�� �� V�����  �����  �  �    ��� �� ��  Q�����"��  �� ��"�� ��"�� ��  �  �� ��  �� �� �����0��$ ��  \������� ��x��� ��d0��!���d�� P�  
���f������` ��*��Y ������  ^� ��`0�� ��	Q���� �� @2  � C� C� C� C�  Q�0����  ������ W�  ` �� 0��p�� 0��0��p��0���� ����� ��`0��!���d�� P�  
����8������ ��3��(�� ����h���0��0��% �  ���� �� ��8 ��� 0�� 0��%���8 ��P��82 � 0��$������P��������@��`��Q��
-��0��@���� ����d����
P�d�   
���l���� V�����	@��|����
P��$������ ��+�� ��� ���0��  ��	Q�	 ��
 ��3�� �� �� �� �� �� �� �� �������� �� �� ��	 ��
 �� �� �� �� �� �� �� �� ��T ���� �� ���� �� ���� �� �� �� �� ��@ �� ��� ���@ �� N� ��  �� ����  W�!$��(��) ��!(��* ��!,��+ ���  ��*��
 �� � �� ��0�� ��g ��. ��o��0����� �� 0�����
���0�������� �����'���0�����
���0�����b���0��
0�� ��� �� ��p��p��p��p��	p��
p��p��p��p��p��p��p��p��p��p��p��!��" �� ��&����# ��+ ��'��n��$ ��; ��(��d��% ��)��*p��+p������� ��!���d�� P�  
��t������ ��*�� ��`��e � �� ��.����� ��0����� �� 0��0����0��0����0��0����0��0����0��0�� �����	��
���� �������� ��������� ��!���d�� P�  
��C��� ��*�� ��`��5 � ��0����0�� ����0������ ��!���d�� P�  
��-��� ��*�� ��`�� � ��0����0�� ����0������ ��!���d�� P�  
0	���� ��*�� ��`��`�� � ��0���� ��0��0����������� ��!���d�� P�  
�	��������,����`��0��  W� �0��$0�� 0��0��3��3�� ��$��� ������\������ ���������?���l`���������o3����� �����$������$���,����]��.Ƞ�.��^���_��3��	3��
3��3��3��3��3��3��3��3��c��m3��n3��   ����*�� �0��  � V� `� �`��� �0��x ��F��F,��  V�F������� ��$���0�� ��!���d�� P�  
�
娿��l���  ^� 
0��3��0��3�� ��m�����P��0�  

P�$�0 �  

P�4�00�  
	P�à0��  
0���	P��0���0 �� 0����3�� ��3 �� ��	Q� ����0���,$��#��,(��#��,,��#�� ��#��������3��3��!��3�� ���3�� �����3��
P�3��B<��3��B4��B(��#�� ��3�� ��0�� �� ��<0��0��@ �� ��40��	0��, ��
 �� 0��0�� ��A��0��y0��( ��B��(0��t ��L��x ��N��H ��< ��@��P ��@ ��@��D ��4 ��@��T ��, ��@��X ��  ��@�� �� ��@�� �� ��| �� ��@�� ��I����I����I���� ��, ��A��� ��( ��A����(���������( ����B��0��B(������#��L$��t ��LȠ���N��4����#��N�����x ��#�� ��8��<�����< �����L�����<���@Ƞ�H ����@���N��(���< ��@ �������P ��@��4�� ��#��AĠ�A(��<��@����H��(�����,��A��4������,��A��D�����	��,��
0��D ��  ��@��@ ������ ��A�� ���#��T ��<0���#��0��H���C4��(0��H���4 �� ���#��0��@��C4��0������X����������,0��L�� ��L0��"Ġ�"��@ ���#�� ��"<��  ���#�� ���#��< ��P ��( ������#�������| ��T ���������� ��� ���#�� ��X �����������3����	  �+�� �� ��\ ��"4���3��"8���3��"<���3��  W��  00����*�� ��#2��00�� �����?0����0�������1���� ��2 ��� �� 0��{0��0��90��3 �� ��0��g0��0��l0��0��0��� ��,4��<"��0��,<�� �� ��0��0������4���� ��5 ������6�������7���� ������8 ��p��p��p��p��p��p��0���p��p�����p��p��p��p������9���� ��: ������;�������<��� ��= �����>������C��@p��?���Ap��Bp���� ��!���d�� P�  
`��<���0�� ��*�� ��0C�0��, ��������� ��
��0�� P��r �����Q�  ��)$�� ��| ��)Ƞ����)̠����0��  
  S��������� ����0����� ��!���d�� P�  
������ ��  P�k  
0�� �� ��*��#5��0��� ����	\�  ����;��#;��  S� � � ��� �� ��`�����0B����0l�����0��:  �  ��F4�� ��*��0��F8�� `��0��F<��0�� ��� � ��8��0�� �� �� ��ʃ����	R��1 �!�^� ����� ��!�� �����!��!�������0��  
 S������ �� ��0������d�� P�  
x���������k�� ����� ��`�� �� ���� �� ��0�� R����������4��a���୽���� �� ����0����d�� P�  
��墽��$������3`��  W� N���� ��r��(��,<��/5�� <��0��0��������?���#<��0�� 0�� ���5�����5�����@��`����������������"��)���"��",��*���+%�� ����,%��,$��,Ƞ�-%�� $��.��� ��0��1%��2�����5��5��e��,��	5��,$��
5��5��e��5��5��5��5��5��5��5�����3��� ��5%��6��4����7��  �� ��h���0�� ������d�� P�  
� ����I���p��\��� W�H���p ����� ����� �����d �����` ��޾�� ��ܾ�� ��ھ��
 ��ؾ�� ��־��  ��5ލ����� �� ��0�� �� ���� ����d�� P�������;���X���o��Æ���0�� 0���0�� P� P�/���� ��@-�@�� ��  P�  
 ��  Q�  
������� 0��0��t@��  ��  P�  
���� 0�� 0��X@�� ��  P�  
���� 0��0��  ��0��80��  ��,@�� ��  P�  
���� 0��0��  ��0��0�� ��  ����� ��8���@-�`��0��PA� @��`��$�M�(��0�� ��c��p��q- �  ��0���� ��0 �  P�  
(�� ���- �`��P��
0��`��S��  U�0��P���S��@�� ����Z- �0����0�� ��f���- �0�� �� ���� �  P� �$Ѝ�����8@-�W����� @P� �8�� �� ��� ��0�� �  P�  
�#��S?� R�  �0�� ����T!���@�� ���0��P�� ��XQ�����  P�  
,0�� �� @��8���  �唼�� ��5��� �� 0�� �� 0��8��� �é����N-� `��  ��0�M����p��0��0�� R� �!���� ��
 ��r��$�� G�0�� ����,0��- ���  �� ��- �0@� !��, �� �� �� P��1��  � U� 0�� ����� @���  �
0��@��C�����  T�������I���0�� S�;  �ܓ��0��  S�	   �ှ��  P� �����  
�3��  ��@��  �夓��0�� T�  
 �� ������#�� 0�� ��0�� ���0��j���  P� ��  d��7��� ���  �@��T���\ �� 0��
�� P�  
43�� �� ��0�� � @P�\0��� ��  ��"���  � 3����0��@��  �0���0�� S�|  �ز��0��  S�   ��?���  P� ��  
�2��  ��@��  �夲��0�� T�  
 �姽��"�� 0�� �� ��0�� ��0��*���  P� ��  p��]  �@��\���` �� 0��
�� P�
  
<2�� �� ��0��B �  P�8�N  
`0��:�� 0�����0��  S�   �����  P� ��  
�1��  ��@�� ��ܱ��0�� T�  
 ��u����!�� 0�� �� ��0����0������  P� ��  ���+  �@��  T� ��0����� ��	��B!��p���0b� ���0��0�� ��I, � �� ��� 0��( �� ��
�� P�  
 �� ��0�� � ���  P�8�  
0��( ��1�������� ��	��, ��0��0��A��  ��嘻��4  �  T�2  � ��, ��0A� U����  $ ����, � �Q�   ���0�� U� @�   ���� - �
�a�@��  Y�  
	 ��
 ����0��� �  P�    �	�� �� d�i �0��P����@d� ��0������ �� �� ��0�� U����� ��   �  ��0Ѝ����� ��͂��8������*���^��Ë��ÿ������,��� �� 0�� ��  Q�  
 ��  P�  
 �����  ���/� ���N-�����M� @��(�, ���00�  Q�  
 ���  �  �� ����L���  P�����  � ��
�� ��$0K����  P�y  � [�  R�q  
0��4��~?� ���M���0��q�ᇑ��	0�����  P�_  ڌ ��J��� `P�[  
  �� 0��$�  ���� [�1�� [� R�  
 R�0��  
 R�  
 R�  �  �� ����� 0P�.  
�0�� �� ��:�	S�  


S�  
	S� p�    �p��  �p��   �p��, �(0�  R�  S  
0 �  R�
  
	 ����9 �  P�#  00�P��, � p�� `��#  �0��  S�    �� ��$����� 0P�0��0�   ��P��u��� ��  � W�t �  
 W�l �  
 W�d �d �ƺ��	 ��\ ����º�� ��c��� ��  �  �� P�� P�4��  �2[����0�� Z�~��: P�� ���K�����#���*���8���1���?����N-�����M�`����� @��(0� �0�� 0�$`�0�� ��0���M� ���@�� �� �� �   �@�� 0��/ S����
  S�$0 � 0�  
 ��/��� � �P�
0�    �  �� C���� ��/ R����
 0� S��$    K��� 0K�p2� ��+���  P�e  
 p�c  
 0� S�Q  �!��0��0��0�� S�  $ ���C��� ����@���  ��R  �$P�0��  S�    �� ����k��� @P�  
 �� �‼�� @P�  
 ��< R�  �,��o �	  �0�� �� ����� 0P�   ��@�����  �0��  �� ��$ ������  T�   ������� ��&  � 0��/ S�   �������0�� p���p����$ K� 0K� ��y��� P�� ��Ż��  U�   �������� ��  � ��������  Z�  
 0��
@��  S���$0� ��( � 0�� 0� 0���K����� ��@-�@��h0��  P� ������  
0������#�R���  P�  
 T�   �� P�  � �  � T� �   �� P�  � �   �  ����� �È���@-� ��  Q�  
 �� �����0���"��������  P�  
0�� ��  R�   ��  ��������  P�  
0��$ �� ��0��  �0�� �� ��������  ����� ��@-�`@�� ��  Q� �  
��� ��0����� P�  
8 �巹�� ��	  � �� �� ��0��g��� �� ��������  ����� ��H���  P��F-��M��M�@�����  ��1���A���� ���Ā� \�  : ���嗹��Q  �Lp��  W�  l�呹�� ��S  �k���T��k��  V�  
 ����� �� ����	0����`�� P�(�9  ,f�
 �� R� ����@b����P�� �  T�7  
���`��p��  W�  L��� �� ��0��p���� ����`��
 ���� �� �$  �L��委�� ��
0��	 ���� ����`��	 P� �  �T�  
 0��L��L��� ��P��0�� �� ����`�� P� P��  
D ��D���  ��  � ����	 ��\ � ��   � ��Ѝ�ۍ�������g��Þ���Ʉ��������@ �� �Q�@-�L ��   �������0��0��  �����  P�  ���0�� ������� 0��  � Q� ��0�� ��AB�  R�  ��q������/�8@-�<@��0��P��  ��  R�  
`�����  \�  
�� �� ��<�/�8���  ��8���l�� 0��  � ��� B�  \� ������0��  R�����/� 0��  �/ R�\ R   `��/�0��  ��  R����  ���/� 0����� ��0�� \�  
  ���/� S����  ���/� <��p@-� S� @��`��
  
  S�  
 S�H    � ����`) �<�� P��  � ����Z) �<�� P��ef�  �U��eA�<�� U�  
< � ����0�� ��0���� Q��#�5 �����  P�(  �\�� <�� S�`�� �p��  S��p�� S�   ��0�� S�&a��  
 S�`�� � �p�� S�0��`� � �� �0� 
� � 
��p���0���`�� ��0��  �#4�� ��p���  ��p��� 0��0@-�@�� ���0��@��@�� ���@�����  \�"  

 S� @����� ��� 0��P��0�� @�����P�� P��@��P��  U�  
 S� @�����0��0�� 0�����  \�
  
0�� 0�� �� �� 0����  Q�0� 0�  �0�� ��0��� 0�� �������3�� �� R�s0��s0����� ���/��@-��M� P��p��@��  ���� ��,���`��  P�*  � ����@ ��W �1�� �� ��  S�1��@P�$P� 0� 0� 0� 0���J � 0��0��`�� 0��  S�  ��P ��;���  P�  
  �@ ����5���  P�0�  
��( ��/���  P�  0�� 0��   �  ��ߍ�����C���L���U���p@-�A��p�M� 0��  S�� �*  
� ����� 0�� 0��0C� S��  �B�� B��(B��0B��8B��@B��� ��
  �� ��  � ��  � ��  � ��  � ��   � ��@�����DP�� �� 0�������  ������ ����l ����� @P�  
t ��ٷ�� ��  �``���� �� ��� �T�� ��0��L �� ��k@��[@��ʷ�� ��pЍ�p���l��^���q��Ün��*[�ån�ën�ïn��~��Å��Í��Ü���@�ô���  Q��D-�P��@��< 
, �0��p�< �p��d���M� ��1'�� �����  P�  ��[��[��  U� �  
 ���� ��������  P�  ������ �� �  ��   �  ��܍������D-�  Q�p��P��
<  @��0�;��@� ��� `��  ��4�	 T�0�� ��  �T  �  T�	  
  �� P��  � P�r@��L   U� D����:J  �@��*  �
 ����� P� ��  � <��  S��?��2� P�  �� ��d���8  �
< �
 ��0��� ��4�����  P�ؠ�  
.  �  �� ��� � R�s@��(    T�0D����
@��   �����0���� �� Z� �J�
 ������ PE��� �� �����  P�   0��@ ����
0��  �� �� 0��� S�  �  
 S�:0� 0� ����� ����  ��J �  ��   �  ������  Q����
����ׅ��t���A-�P�� `�� �� �� ��: �@�� 0��0��   �@�� p��  W�  W p�p����0��  S�  S  
.0����0�� �� ��% �p��   �@�� 0��  S�  S���  ��  �� 0��� S�  �  
 S�:0� 0� ���A�������N-�Z�M�0�M� @��Y��P��(��Z�� �� �����.�����00��  P�8 0,����  R�p���̍�, , ��������̍��,��00��T ����, 㲠��Q ��*�0��  P� ���
 � ��A�z���̍������V ����"U���"  �!"� � �� 0��@<��   �@�� ���/ Y�\ Y �������
1m����`�� ���
 � �����D|��  W�    U��g�P�� 
  � �����  P�  �Z��0�� 0�� �� `��l�C�   �`�� 0��/ S�\ S���
p��  �  U�g��p� p��?�p��p�� ��������������� `��0<�� ��  S�`'���>�
0����e���  P�� �DG��p  � �T�,�� 0��� [�D0��g  
0T� �  
 �b  
@ �`  
0��0 �����
0��  Q��&��U}��`T� ��p���� p������ U�  0T� �̍D0�(  
  �  [�   U� ����� ����J��� � U�  
 ������ P� `��;  
`��Z}��
 �� p������� U�   T��� �0��	  
  S�,  
0����/ ��0��0��0��,���$  �  S�"  
��� ��� 0����������!���  �1�������� ��l
 �  P�  
U�� ����f
 �  P�  p�� `��  W�  
0�� �` 
p����������  �`�� @��p��%�� �D� T���0<��  S�  �N�����
@��0�� Y�
  ��0 ������>��0�� �� ����0�� ��0#�  �0��0��0��e��� ��U͍���� �� �� �� ������  P�  ��  ���� 0��
��� 0��   ���� 0��/ S�\ S���
  Y�  
���  S� �����
  �p��  Y� p�p  W�����  
 �������p��  �� ��0<��Z͍�0��� ���  S�`4��Z����X$�0��0�� P�,���P��/�p��$ ��X�P���>��0 ��
0���� $��0��4������ �P�  D��i  � 0T�ˍ�  ��� S�D ��a  
 T� �  
 �\  
@ �Z  
�T����#��Q}��0��p��$��� p��������  Q�  
0T� �+�D0�(  
!  � 0T�  S�	  ��	P��p��  Q�\  
�� ��D��t���W  � ��  R�  
 �����$0�� P�3  
Z}�� �� p����B������  \�  
0T� ���0�  
��/ ��������Y���   �  S�  
��� ��� 0����������N���  ��� ��	 �  P�  
Q�� ����	 �  P�
  U���� ��  ��,���p��Y
 � ��  Q�*  �$  ���� @���>��  D�
0�� ��0 ��0��Z���:��O��� P� P��  �0<��  S��?��2� P�v��:��	P��p�����  �p��	P��0w� 0�3  U� 0�  S�P�� ��h  f  �̍�O0�� �b  

`��U������  W� ��0 ��
< ��� ��㳰��0<��!��  S�0�勴��q�@��(���x�  Q� Sp��p������  � �������
 ��0�� P���E� \� ��"   U�@��<  �0<��  S��?��2� U�6  *p�� ����0`�� T����:@k��� ��
 ��0�����  P�  0�� ���� ���d�0�����  P�	�� ��   

  ��������������d������@��  P� ��  
� �庴��  ����� P� P�� ��  �0<��  S��?��2� P����:D �嬴��   � ���	 ��kލ�ڍ�����a2��t�Ô��
���������Ô�î�������t�Ô��ׅ��#���p@-� @��P��  ����`�ᒴ�� ���� �� 0��p@�����:��� ��0�� �����`����@-�  \��M� @��P��<  
�p��`�� �� �� ��0�� @��<�/� P�  
��� ��s���.  �2��U S�+  2�� S�(   ����/�����  P�2�0��0� P�  
6 ���� �� �  P�  
R ��t�� �� �  P�  X0�� ��  ��  ��@0�� ��  ��� ��@ ��K���  ���4 ��"��2��E���  ��   �  ��ߍ�����l���~��@���p���p��F���V��`����N-�  \��M� `�����  
�E��P�� �� �� ��0�� `��<�/� P� p��  
��p��$��� p��F �
2��U S�  2�� S�  
L���  � ����/�����  P�2�0�,5� ��  
6 �� �� ��i �  P�5� � p�  
�� ��������������"��2�����������)��� PP����  
 ��,��� � @���� �� ��0����@����d�� P���    T����p����	 ��0�� ��� 0�� ��m0��0��o0��0������0��  ��`�� ��0��0��Գ��"��0��R�D�5�  :R�  �8��
���ʳ�����  �R�  � �����0��³��0��  �R�  ��弳��0�����0��  ��R�  ���崳��0������}R�  ���害��0�����������ᩳ��@�� ���女�� @��0��@��0��  ��@���� �� ��@��$���
 ��@��	@��@��@��@��@��@��@��@��@��@��@��"�� ��"Ġ� �����"Ƞ�",����� ��0��$ �$ �� �� $�� ��� �� (�� �� ,���� ��w���0��@��@��@��G ��0�� ��@��30��@�����@�����)���	@��
@��@��@��@�����0��0��@��@��@@����[���R ���� ��W���U0��U����1������ ��0�� ������d�� P� ���r  
X��I���#���P��������,��: � p���A��A ��r��������U0�� ��U����1�� ������R0���!��a���0��
 �� 0��0�������������q���q���q���q���A���A���� ������d�� P��K  
A  �h��?  ���,�� �
��E��� �P��7  
��*�� 뉐��|��  ��� �� ������d�� P�\��   
��� ����$ �@��  Q�  <������	�� �� Q�
0������$�� p��������p��0��p�� �� 0��0������p��p��p����p��	p��
p���� �� ����d�� P�  
� ��۲�� ��ߍ���������� PP������������� PP��������� ��˲�� p������l���~����@���p��F���V�Ä��q��Ô��Ü��ï���؆���������������������*���;����p��D���[��À��ã�������ч�È��Ëd��������0��  P�  � ��/�8��È��� 0��p@-�`�� @���M�P�� t�  h �嘲�� ��  �  ��/ R�\ R  �  
 ��D�� ��@�� � ��(0������� �� 0���0���������ۍ�p���D��#���J���,���x ��0@-��M� P���M� u�  ` ��r��� ��  � 0��/ S�\ S  
 0�� ��<�� �� �@�� �� 0����$ �� 0��##�����Ѝ�ۍ�0���D��P���J���,���8@-�4@�� 0�� 0��,0���� �� PP�   ����h � P��0��  ��8���D��,��á��@-� 0�� ��/ S�\ S�1�
     ��� 0��/ S�\ S���
�! ���X �i  �0��  ��  R���� s�/ R�\ R  � ����
@��  ���  ��� ��  ��. P����
  P�  
\ P�/ P  
  ���  ��@��/ P�\ P���
 ���. \����
  �0C�  ��\ P�/ P�����  S�  1��
  �0C�  ��/ P�\ P���
 B�  ���  ��  R����  \� ��� ��  �0��  R� �/�� 0�� 0��%  ���� �� `�/ �� ��0��  �0�� ���! � P�  ��  ��  �  ��  ��  ��  R�   S�  
S�/ Q�\ Q C  �/ R�\ R  
  ���  ��/ R�\ R���
����������  �����H��I��G��D�� 0��@-� ��  �@�� �� ���#D$��@�����4,�s0�� R����� �����D���0��@-�0�  R� 0�0P��  S�
  
��� R�0��� ����1�� #�  
 ����P��"��`E� � @�����  �p��@��  ��p �q�� '��p �q�� '��p �q�� '��p �1�� #�  \�80���L����  R�1�������� R���0��� ������ !��������D���@-�  ������  ����������N-� ��������� P��<@�� ��
 ����# ���  
�p��`��  V�    �
 T�P��
@D����
 ��0��| �� ���W���Ѝ����� �� �� ��# �  �� 0��  ��
 ��0��
 �0�����
@DP� ��`��" � ��  ��@�����	 �� ��Ѝ��N��:���D���x��Å��É���@-��� ��2���  �����\���	���N-�P�M�p��P��p@�� �������@ S�  �@ ����! � @��  T�>   ����! � @��9  �� ���� T�@�!���	��� `��  � U�0�  �!�  
 U�0�� �  �� � �� �������`����� V������:�� `�����
  � ������ �  
� �  
 ��.����`�� V������P ��P ��0��  ��D C���낱��  P�  �  ���pd�  �0��0��  W���� ��PЍ�����3�Ñ���H�×����L-��@�� p��`�� Q� ��� ���  � �� ���\! �
 �� � ���@T�P�� �� 0�� �� ��  � ��0��  ����  S� `�����  �    R�   
`�� U�  �   T�   ������� ���� S�  �   R�  �@T�P�� ��������` �����  
�0��b ��������� �����������F-�D�M�@�� `��$���p����������P�� �� ��<0��(���d��� � P�  
� �傰��  � 0���� ��p��0j�`��0��
������ �`p��0P�0� W� �� 0�  S�p��  
@ ��l��� �� �  ��  �0�� ��`f� `�� � ��DЍ�����Da��<a�ß��å���Ȉ�����7@-� \����  � �  
� ��  � �
��
��@���Č �  
@��P�����  U���� �  
@��P�����  U���� � ����� \�  :  ��#���  ��  ������� ������>���������� ��ϱ��� �� ��V����@-� @P�P�`�  T0�� ��  ������ 0��p��0��P��  S�  
 �庱�� �帱��0�� V�`������  �岱�� 0�� 0������t��  ������x��p@-� `Q� ��0� �  
 0��  S�@� 0�     �@��P��   �P����� �� S�  *�  �  Q������ ���  �  Q����
 0��@��0�� ������� 0P�0�  �� ��p���t�� ������x���N-�����M�  R�$ � P�� � ��p��!�� �� ���M�@�� `��� ���*    �� ��7  � ��0����  Q�   
 ����, ������(0�3 � �(0�  Q�, � ��� � 0�   ��) �, � ���
  � ����� Q�  
\ Q�   �����0��  Q����`����� �����0�� R����� ���� �� 1��i ����  W�
p�  

 W�  *  �� ���0��  ��:  �$� P��  U�  
 �� �� ��y � 0�� ��*  � ���ჳ��$0�  P�  �� P����������  �� ���   �E� ����� ��P��  Q����
P��= �� �� �����	  � ��
 P�  
\ P�  \ �� �� ���� �� ��  P���� �� ��0����� R����� �� 0�� 0���K������d��t�����0�� �� ��  ��i���x��  �� 0��  �� �� ��N-����P�� ��� �� ��0@����� � ��� 0��  � s��J� ��  Z������:  � �� 0��  Q�`�`��� ��0��  S�p�b  
 S�$  �� �� 0��l � 0��  P�   �� R�    Y�  
  �� �� �岰��	 �� `�� �  ��`�� 0�� �� �� ��  R�
 � ���1� �m  
  �� ��p��p�� p��h  ��� ��p��A�  �0�� W�pc� �� c�p�� �� W�
�,  
  ���� �� R�#  �� �� 0��3 � 0��  P�  0�� S�    Y�  
 0��
0�� ��y���	 �� `��` � 0��`��
0�� ��0��  S� � 0� ��0�5  
 0�� �������� ���0  �  ��
 ��  R����0�� S�#   ��0�� R�  
0��  ��� �����`��= � `��`�� ��	 ��8 � 0��p��0��  S� ��  
0��  S�    �� ��  ��
  �0��p�� ��0�� p��0��  � 0�� �� �� 0��0��  ��Ѝ�����t��0@-��M�0��@�� ��  �� ��0�� @��D��� PP�P0� � �  �  
0��  �����0�� �����0��� 0��  �� �� ��0��0C�0��Ѝ�0���t�� ������x���N-� `P���� �M�@��p�� � �  
	 �ጰ�� �P�  
 �� ��2��  ��~  ���	 ��r �@0�� �   0��  S�  
 ��#��� 0��  S�  

@��  �����@ ��P���8��� @P����
 ����� ��b  �@�� 0��  S�	 SP����
# S�0�	     �@�� 0��  S�  
 S����P��G  �0��  ��  R�= R  
 R����  �  R�P�  
��P�����  Q�  
 R�  
 Q�	  = R�P� 0�0� 0�� ��0����}���)  �  ��P��  ��0��	  �\ R�  �� ��  Q�    ��P�� �� ��  ��  R�  
 R������  ��  ��0��@�� ����� �� `�����0��  S�  �� ��D ��0�����0�� ��	  �P��	0�� U�  * 0��  S���
 ��|��� �� Ѝ�����t��$���@-������ 0�� �� ��0�� ��a������x��@-����0�� �� ����� ������ ��Ѝ� ���x���/� �� R� ��/ �� P�  �  ��/�  ��0��@-� B�1��  ��@��� Q�0�������:  ����� 0�� ��T0��P ��0��0�� ��X0��\0���/� ����N-� \� @��p��P��   ��  P� ��f  
���@�� `��@��  ���������� [� Y	 ��0��  �X  
����0��  P�	  �@�� ��	e����1����� �� �� ��  �  
@��������1�����  �`�� V� �������:@�� ��� ���K��� V�  *��� ��1��0����1�����`�����!��0�������������  P�  
0��`�� ��
��`����� ��  �  Y� �   [�  ��  ����0�勱��
  � ;� W��50C2 �5�50�"�!� �q�'P�%  *  S�����0��  �� W� 0��p�50��P�5 0��Ѝ�������� 0������D-��� @��Pp��P��`��  �X`��\P�� ��P�� Q� V�  �0�� S����: S�  ���� V� `�`� U� p�p���P ��  
��O���  ������  V�  
0��
 ��������0�� b� ������  W�0��  
�A�� ��0�� b� ������!��A���b� a�����D��L���P ��J���p@-� 0�� @��  ��  ����`��0��`�� Q�  * \�  *p��� P�P�����:  ��p��� ������ a�  ��/��N-� ���P��P �� ��@�������� B�  �务��4  � �p� P�,  :  [� � �  d   
 W�%  * ����  [� d�  d�  �������  P� ��	  �@D�  e�P��	 �� ���	���  P�  �  �0���� P�  d�  :���� �� `�� W� 0��0��  V� ��	 �� 0�  S���� 0���J�0C� 0�� 0��  S����� `�� ������0@-� 0��P���  ��  �X ��\@��0��@��@D� Q� P��P��  Q� P�3  U�  
 ��0��� R� �����:  ��0����/��/�p@-�P��@����� `P�  �� �� ��b��� ��p���U��� 0�������@-�@�� P���� ��p��l ��� `�� ��� �  T�  �  Q�g�`���� �� `������s@-� @P� �  
 `��P��  T� ����
 ��   
 �  T��  �`��T��  
@�� 0��  S�@� V�������L�%���X���%��|����N-�  R� Q�M�`��@�� ��0��=  � A��� � P��0���P��  U����:����`����0�� ��� �������� 0e� ��	`�� ��p��0��	 �� ���
��� �� ��0�������<�/� ��0��  P�  � �� �������� ���� T�������p�� y�`�����:�����0d���� S�������: d���y � PP����Ѝ����� 0�� ��  R� ��0������/� 0��  R� B��/���  \����0������/�  ��   � �� 0��  S�������  \����0������/�  R�0@-� 0�  0���0�� ���  \����  � R�    ��  ��0���P��@��0��  T�@��������0��� 0����� ��0�� b�r ��  R�    \����r ���/�@-� 0��	  �@�� B����0���l�|���  \�    T�  
  R�������| �����  �  S� ��   ���/� 0��q �� S�����/� 0��   �0��  ��  R���� `��/�8@-� @��P������  ��  ��u0�� R�8�� @� P����*  ��8��� 0�� Q�  ��  
���0��  \���� `��/� 0��  ��@-�  � \�  
@�� ��  T������� �� ���  \���  ������  � S��/��� ��  \���� �� 0��  S�  ���� ���/�8@-� @P�P��  `0�� @��  T�  
 �������� 0��  S�< �@� 0�
  
�� ������  P�  
 0��  S� 0�0�0��  �� ��8�����8@-� @�� P��  T�  
 ������  P� 0�0�  �� ��8���  P��/ 0��  S� � 0�  �/� C�C� ��  Q��/ ��0��  R�����/�0� ���@-�  @��0����� S�D�������� 0��  �@��0�� \��L�������� ���� 0��  ���0��  R� B������� 0��  ��  � ��� ��� �� R����* ���/� 0�����0�@-��� @��  
	  �@��@��0�� \��L�����@�� ����@�� 0��  �����0��  R� B������� P�@-� 0��  �  �������0��  R� B������������ 0��  �@��@��  R�0C� B�������@-� 0�� ���  �@�� B� �����  T���  R���� �����@-� 0�� ���  �@����� T��� R� ���������@-� @�� ��p��
��� `P�  
 ����� P��  �����  P�  
@�� U� ���� ��PE����� @�� ������  � ��� B� \��/ ��  R�q0����� ���/�8@-� PP�@�  
���� �♬�� @P�  
����� ��8����@-�}_�� @��H�� ��u �@�� `�� �� �� ���� p��( ��V �k �  P�  
 ���� � ������@B ������������8@-� @��P�� T�P�1 ��gx��@T����8��耖� 0�� 0�� �  @p ��/�H��0����  �����!2��0�� ������/�L����@-� 0�� @��P��0 S�`��  0��x S�   ��0���� ��D �@�`�    V�`�  �  R�
`� p��  �7'�@��  ��@ ��00@�  ��D �  
 �   �70@�  
����70@� S����:  U� �� @�����H��@-� ���- \�   ������  `����@������@-�@������ 0��  ��K R�
  
  �G R���  �M R�  
k R���  � �� �� �� ��i R����� ��B Q�  �0� 0�����D-� 0�� @��P��0 S����  0��x S�   ��0���� ��D �@���    Z���  �  R�
�� `�� p��  �7#�`��@��p��  ��X ��00@�  ��D �  
 �   �70@�  
n���70@� �����  Q�    Z�*������  U��� @� ������H�� 0��  �
�� ���##�  �����  ��0 B�r��	 Q����� ���/��D-�Q"��QD��!6�����P���`���������Q!�	P��#%�
 �� p����T%�e��P���a�0��������� ����@���Qe���0P��P����������Ad�1��0@��@�������Š�  \�<c�0��00��0�������� -�@-� ������N���
 �����  �����  �� ��  �� 0���y��@��Ѝ��/᠆ p@-�  Q�`�� @��`���P�� ������0�� �0�  ��  
  � ��C�PE�@����0�� R����� 0��  �����0�� S�������0��  � ��C� R� ��PE�0������p��蔉���@-� @��� ��p�� �����  W� `��  �0�� �� V�  � �����������  � ��P���� � ��  �6��� P��U��U2��%�� ������ �P��	��,%�� ��1.����
0�����.�e������Ve���0P�� P��P��Š� ����l�� �0������à����`���0 �� ��%��0 �� ��a�0����@����꠆ �� �N-�X�M� @��P��x��� �|`��
�Y��� �%��P� ���  
  S�  � �  
  �  r� 0��`F�-p��  �`F�+p��  � �`F p�    p��  [�  
 Y�`F�`F��00���0�  

 Y�  
 Y� ���I�������������P1�� ������� ��|0��0�����0��
������B �  ��0�������  ����
 ��o��� �j��0�� Z�
0��0�� �`c� �  
  � ��B�`V�@�� �����Z  W�p�  [�  
 Y�0 �� ���X � � �   � ��0� �   �B�`V�@�� �����Z  �0 �� D�0C� �� Z�@������X0��
��EA�  �0��0B��Z�0��A� �����Z  �  �� C�`V� ��0�����ZXЍ�����L����N-�P�M���� ��� ����r �% S�.  @��0�� �� ��0��+ S�  
  �  S�  
# S�  
  �- S�  
0 S�
    �@������@������@������@@������@������0C�q��	 Q�  � ��
P����� `��
  �* S�
P� `�   `��P�� �� ��  V� `f�@��0��  ��. R��� p�   �� ��0��0C�q��	 Q�  � ��h��� p��  �* S�   p��P�� �� ��  W����  ���� p��0��  ��h R�l R  
L R�  
Z R�  
z R�  
t R�  �  l R�����  0��l S���L ��� 0��n S��  
  �c S�  
  �% S��  
X S��  �  �d S��  
i S��  �  �s S�!  
  �o S�  
p S�  #  �u S��  
x S�  �  � �	0�  
  �  �� C�`F����  V�0������  ��	0�� ��  �  �� C�`F����  V�0�����ʍ  � @��	 �� �� ��0�����Y����  �  ��  R�	 � �0�H�%  
0����M S�  
  �I S�b  "  �i S�  
m S�]  @@��$�� ������ ��
��T���@0$�S3�� Z� 0�0���  S�:0�0� Z���� �� ��	 ��0�� ��� ���$��@@�� @��)��� ���M  �@@��0��6 S�  $����� ��� �� ��3�����1���@0$�S3����� [� 0�0���  S�:0�0� [��������4 S�@@�#  $���0�� ���p�� ��LP���� �� ��0����� �� ��0��  e� ���  ��|������ \���� [� ������.�� [����P�� ��p��	 �� �� ����� v�	 �� 0�� ��	`�!�`������p�� ��K��������0��`!����0��0�� �������D  � �����	0b�  �� 0��>  �0��<  ���  � @����  �@��  �%0��0��0��  ��  R�0C �0�,  �
��L R�P�P���� �   
l R�    �� ���� 0��  
  �Z R�z R��  � 0�  
t R���  �  
h R����  ��0�  r ��  S� 0��r �    �  S� 0��   
�?��	 ��� ��@������ ���0��0��0��0�� 0��  S��� 0��0��	 c�PЍ����蛉��H�� -�@-��� �� ��t���@��Ѝ��/� ���N-�`��T���@�M�LF�X���`a� ���(��P��p�����0��Y���L�pG�0C�@D�p��`��@��PE�$���K�,p��<`��,p��(@��4���4P��P`��LP��0���8@��<��8p�� ���0���P��`�� �� �� Q�  � ��P����� �� ��A����B��4p����� ���Q��	p�� �� ��  U�4B��b�  ��%�� ��  
  �� �a���  
P�  ��  
 Q� �5A�0  ��%���2e�4E�� �� Q�  �P��`����� ��P��A����@��0P��`�� ���� Q�� a��p�� �� �4@��`�  ����  
`� Q�  * ��A���� Q� �5A�0�2<��� P��V��f� i�P��  U�4F��`  �8`�� `� P�  � ��P�� �� P���R��  � ���  Z�pI�  $��� P�	``�p��	  *`�� ��� ��� ���[� �����	0�� i�pe� ��5  �  Z�   *$��� `j� V�	����`����p�!���* f� �����0��0��`�� P�0��`��0�����0�� Z�	0�����*`�� ��� p�� ��  Z�p�����
0�� j����� P�
``�p�����*`�� ��� ��� ���[� ���������0�� B�0��0��0��0��0�� R� 0������  R�M  
 �� R�p�� �� �(  
F  � � e� B`�`� U�pC�  ��P��`@�`��`�����`V���� ����᱐��0������0��p�� �� ��
  � U�PSᢐ���`�%T�	`��`V�P��0������0�� �0��  
 �� ��  �p��@ �Q��a� ��p�T��
 ��P�� �� P��P��P��  �@ �Q�� � ���
 ��  � ��P� P�
  P�� P��|P������(���, ��	 S�  \1���: �� ��(p��a��,����f�\��A�P��p��Pc�P�� P��pl�A��p�����0��<��8@�� ���0��@Ѝ����袉������։���N-��M�@��0�� 0��0��h�� P��P��0��  S���� 0��  �0`��p�������Q�����A� S���0�����:������ ��删��0��2S�  S�  
  Q�0�    �Q���������@��� @��  ��  ��0������������P��@�� ��@��  �� �� �`��P��RU�  U�  0�� S����h`��P�����p�Რ��p��Pz�	 J	 W����  U�  
Pp� P�3 Q�P�  U��  HP�� p��t��p�Ⲡ�Ა��
��ഠ��P�� U���� P��
  �0��删��p��  W�p��dW����G�`��P�P�� U�`�����:  P�  
 P�    ����@��$@�� ���  �x#��\�� P��@`��$`�� ��  �`s�� ��� ���@���$���p�� Q���1��� S���!`�� P�  � �l��< ��[V�  �3  " ���  P� F�8 �����  @�� ��P�� 0��@��(0�� 0��  ���� �����������pc� ���wp��4p�尠��	 Z� ������  �$��Ŋp����� ���`p��p�շ���p��p�����pc�w�����,��� �g�@������	�0��D���,���0���	�g��g�������������@0�岠�����40��������  \�0��D���0��0�����pB����	���0��w��   �p��  ����  W㈐���G  
 � ��p�ఢW��J�z���  Z�p�   R�Y  
���0���p��p��p�ሰ�� W� �ఢB����8���(���	  �
 R���
  S����h���0�@c�������0�劐��������  �0������l�  [�0�勰��  �@�� Z�������:���	���d��<���0��[V� ��3�
"  Z�5  ,������	Q������k�A�����I���( �岐��v���  S�  
8@��(p�� � Q�|��P� � 0�0C��@���pB������@�� ���w����岐��   �p��  ����  W� �  
G�  � ��   �4���  P����������� ���a����� `��  �  ��   � ��Ѝ�����n������� P�@-�  
0��  S�  
  ��S΃� ��@�� �� ��4@��I�� �� ��L���@��  �� �� ��  ��( ��, ��0 ��8 ��< ��l���P������ �����  R�p@-� @��P��5  
  ��1 R�< S  � �/    P�%  
 0���� ��0%�  S�(0��0� 0�$0��  S�0�$0�( ���� �� P� �p��  U��� Pe� 0��0��  �/ U�E2��P�0��0��0E� S�  �( ��  ����$�� 0��0�� ��p��� 0��$P�� ��40��p@����� ��p���`���X���0�� �������@-� @P�  
 ��  R�  
$0��  S�  
4��  Q�  
( ��  ��3�/�( ��  ������$��  �� ����� ������@-� R� H��`��p�� X��$H��   0��@���?� T��?��LD��@D�P�� U��\E��PE�������  Q� ���� R� 0��  �P  � ��0��@��P��  V�`F�����?� T��LD� �����@D�� �������0��[! � �� R� ��@����  ��P������� P��������P�� �����P����  ��P������� P��������P��	 �����P��
��  ��P������� P��������P�� �������P��  ��@��P���� P��@��P��0��P����� ����P � ��V}��VmF�0p��0`F�@����H �P��5� V����  V�0�� �0  G  �R� R�@��R�  ��P���R��� P���R����P�� R����P��
R�  ��P��	�R��� P���R����P�� R����P��R�  ��P���R��� P���R����P�� R����P��R�  ��P��@R��� P��@��P��P�� V� ��`F����� ��0�p��  ��  ��� ��@��P��  S�0C���� ����� � ��@����� �P�������� �ሤ�� �����N-� �P�`�M�P��� 
@��  T�� 
 0��  S�  0��  S� ��S�� 0��p �����l��� S�D��0� ��� 0�/��0��8`��<P��Dp��4 ��T ��L ��X �� 0�� 0��<���H ��8��T ��(���0�� 0�� S�񟗞 �ė�ü���Й��X���ܚ��|���@������ð��ô��Ü����������ȟ��<��ì���,���,�����Ð�������l������Ü���ĩ�ü��Ô���@��à���������� � �� ��} �	0��@ �	0�� �	0��^  � ��  R�	0�0�  w �  W�� 
S�pG�e��P�� U����0������� ��;� V�  �   R�  
  �� ��  �� P������0��\�� ��`�� ��\0��t0��]0�� ������0�� 0�� ����� 0�� ��  S�  �0 �0�� �  
���� �� ��&��b � 0Q�  
0�� 0��H?�� � � R�%  &b��$ �� � ��  R�0��PE� 0��?��� ���� ��"�� �� ��P������`��	0�0� ��4 ��$ �  W� 
 S�pG�e��P�� U����0�������0�`�� S�  
0�� 0��>��j �
�0� 0��>�e  0��  S�V$�  �0���  
\`��\��&d�� ��]`�� ����� �� P��0��`�� 0��	0��  �  W�Y 
 S�pG�e��P�� U����0������ 0��  S�`�0���  
\`��&<��\��_0�� ��&4��&h��]0��^`�� ��t��� �� P��0��`�� 0��	0��  �  W�7 
 S�pG�e��P�� U����0������ 0��  S��  �&$� �0���  
\`��\��&d�� ��]`�� ��S��� �� P��0��`�� 0�� ��+�	0�    �  W� 
 S�pG�e��P�� U����0������ 0��@`��  S�`�0��<�`�P�  
\`��\��&d�� ��]`�� `�� ��P��-��� ��  � 0��  S� �0�� 0��0���)  
@ ��  W�0�1 0�!  S�   
  ��  R�  
��  Q�  
��� �� `�0�� ��� \� `�  �� ��	�����0�� ���  
 �� ��	��0�����0�� ��@ ��pc����0c�@0��@0��  S��  0��@0��0�� 0�� ��+�$  
  W� 
 0��  �����0��  R�  
 ��  P�  
 ��@ �� R�����7@�5  \� S���: ���  
 �� ��	��0������������0�� ��  \����pc�  
� � 0��  S� � 0��@0��0�� 0�� ��*�$  
  W� 
 0��  �����0��  R�  
$ ��  P�  
(��@ �� R�����7@�5  \� S���: ���  
 �� ��	��0�����������0�� ��  \����pc�  
j � 0��  S�$ �0�� 0�� ���	0�    �  W�^ 
S�pG�e��P�� U����0�������1�� V�0� 0�:�E  P��`�� 0��  �� ��  S��$�, � �0 �  ��x��� ��4 �� �  W�? 
 S�pG�e��P�� U����0������&��&4�����,��<� `��0��P��4��0��40��
0�� 0��0��  S�	    ����p�������<P�� �� ���8`�� �  �� ��  �����0�� 0�� ��4 ��P0�� S� 
0��  S�	0�
  
0�P��6c��0�� �  W� 
 S�pG�e��P�� U����0������� ��`�0�`�� S�  
 S�  
 S�0�  �8��	��T����X����L0��P���� ��  �0�� 0��  �0�� 0��`8��0��"a��PE����� �	0��6b��P��  �  W�� 
 S�pG�e��P�� U����0������8���/�&("�#8�� S�0� 0��7��  P��@0��`��0�� 0��@0��  S� 
 [�0�1 S�0�!  S� 
 ��	��  ��pc�0��}���0��@ �� ������ c��c����@ �� ������  W� 
 S�pG�e��P�� U����0������0� �<�����0��V%��  S��� ��`0��\ ��&g��d��PE�  � Q�  �0�� 0��7�� � 0��h0��0�� 0��\ ��  �  W� 
 Q�pG�e��P�� U��������������PE�a�� ��0��&��h0��0��0����h0�� S�&�%� �   *	������R�0��  ������ S� ������4��  ��4 ��H���h0��0��l��T0��L �� �� ���8���L��<0��������  P� ��0� 0�6�?  ��0�� 0��h ��d ��`0��0��$0��{  �T0��  ��L���	 ��3��,0��,0����� � ��0�� �� S�  �  W� ��0 
0R�pG�e��P������ P�  �  �  W�& 
�R�pG�e��P�� U���� �����:� ��Pc���6c��h����Q  � P�    �  W� 
 R�pG�e��P�� �����  U� �����:  Q�Pc�6c��3  
� ��0�0��&a��&��PE�(  � P�    �  W�� 
 R�pG�e��P�� �����  U� �����:6c�� �� c�0�P��0��a��  �  W�� 
 R�pG�e��P�� �����  U� �����:6c�� �� c�0�P��0��c��  ��$����� Q�  �0�� 0��$4��0��
  �h��0S� ��h ����'�����h��$ ��  Q���: 0�� S���
4��	0��H �� ��8���l��T0��L��<0����L��` ������  P� ��0� 0��3�� l �� ��`��0��8���P ��8��T ��X0��@!�<0����d ������  P� ��0� 0�0� 0�L3�� 1 � W� [�  �  ��
 �����p�� ���8`��<P��(�� ��o���0����� ��� 0��p��8`��<P��q���T0��  ��L��	���3��00��0 ����� 0���1�� �� �� R�$ ��, ��  �  W����k 
0\�pG�e��P������, ��  S�0 ��  
� �  0��  ����@ ��@ �������� 0�0 ��32����1��0��0�� ��$0��, �� �� P�  �  W�J 
0\�pG�e��P������0��Pb�6b��, ��  S�$���0�Pl�@ ��6l���  
  �  
0���  �@ �0� 0��1�& 0�H0��0�� 0��H0��  S�	 �    �  W�& 
R�pG�e��P�� U���� �����:H �� ��3��@��Pb�6b��0��@0��0�� 0��X0��  ��P��	���3��00��0 �����0���!��0�� �� S�$0��, ��  �  W����  
0\�pG�e��P������, ��� �0 ��   ��  ����@ ��@ ��������  �0 ��2#����!�� �� �� ��$ ��, �� �� P�  �  W��  
 \�pG�e��P������ ��Pc�6c��$0��@ �Pc�6c��  
0�� 0��@0���  ����$���	���8���Q���p���e���x��Õ���p�����ù���Ҋ��������։�����â������3���,��� �0��H �� 0��D���H0��  S�	 �    �  W�  
R�pG�e��P�� U���� �����:H �� ��3��D��Pb�6b��0��D0��,0��( ��D ��0��0k� R�0�� 0��0�� 0���0��  �  [�  
( ��D��0k� Q� ���@0��a�  �0 ��0c�4 �� S�0b�c�(��@ ��c� �� S�0�! S�0�!@ ���c�  ��  c�@ �� �� ��� �� �� S����@ ����� ���  R�]��  �  [�h  
  ���K�@0��0��  ��0�� 0��R���0��  S�	0�  6  �  W�Y  
 S�pG�e��P�� U����0������(��0�� k�0��  R�0��0��0��0��  
0�� b�  S�  
 0�� ����s���  � ��� ����?��� ��4 ��0��  S�&$�&��,� �< � 0�4�  �� S�(�� P�`�0�(�� 0�h2  0�� 0��0��  S�  
0��  S�  
	0��  �  W�  
 S�pG�e��P�� U����0������0�� V�  
0�� 0���2�0������ P��`��0�� �� 0�� ��  ��������p��(0��  ��  S� ���8`�� ��<P��   0�� S�L  �0��(��� \�H  
P��40��  S�	  0��$��( �� ������ ��  P�4 ��6  
(0��  S�  $ ����,0��"��00��( ��p��( ��( �� pg��� W�  :b�4 �����  ��(0��0 ��  �00��g�4 ��`c� W�`�1  �� �����pW�  
�� ��4 ��g�����(0��0p��,0��  �00��( ��0��00�� S�,0��( ��0p� S�`�0,`�5  �0���� 0��8  �D ��P��`��(���Pe���0��`f� ����0����0��  V�  R0��0��0��  
 �� 0f���  R�  
�� �� �����  ��� �� ����� ��4 �� �� R�<��P �� �  �  S�@0� 0�P��0��0��,0�� �� P��  Q�  
��  Q����  � �� �� ��`Ѝ����� 4�� ��p ���/��, � ���8 � ����#���/� R�0��@-�@�� ��  �0�� ������0D� ����辋�� �����@-� �� �� ����� �����D Q�C R�F-� @�����  � S�  � 0�� C�r �� S� R  � S�  0�� S�  0�� S�   ������x2�� 0�� P�  
�  ���d������`2��lP�� ��X�� �������� ��A���  P�  
��8�� ��m �,�� 0��  S�  
 �哕��� ������2�� P��@�	�� Z  T  �  S�`�P  
 ��`��`��	 V�K  ��1�� P��P�� 0�� S�  
  � S�  
 S�  
 S�>    � S�'  
( S�,  
 S�7    �1�� 0��  S����0    �x��   �t�� 0��  S�)  �����&  �\q�� 0��  S� �P�     � R�  � ��i���  � R�   ��h���1�� ��  �q�� 0��  S�@��    �q�� 0��  S�  � �� ��^����� ��� ��
 ��~���
P��@��	 T�  * 0��� S���  �� ��j � ����� 0P�  
 0��n S�0� �  �  
������  P�  J	 �  �T �
  �P��t ����F��� ����C���0��  S�i��
e���������p3����� 4��4���	��c�Sc�3��������x3�Ü3�����ü3�� ���|3��
�����ä��#��ü��@-��� 0�� ��0!�;�������N-��q���A�������� �����ȡ��	������� P�����% � �����+�� ����c ��� P�� ��`�������������j����� �p ������ ��( ������, ������0 ������4 ������
�� ��8 ����� ��0�� �� �B��	���c���	 �� ��	 ������} ��	��S �� �� ��	��	0����� ����� �� ��.������	������-������ ���� 0��Q0�� �������0�� ������������� ����i��
 ������� ��  ��  ������ 0��C �� �� ��`c�D0��A� �`�� ���� �8�� � �0 ��: �  ����Ѝ��N��B ������'������L��4�Ä���4���00��@-�0�� S�  �  �偛��@��/ ���� �@��q�����;��Ä��� 0�� �  ��/�� ����� ����0�� ��0��0�� ��  � ��/�  ���/�0��  ���/���80����  Q�	  
0��  ��  R� ��   ���/�40�� S����  ���/���@ ��0��  S�  ��/  ��  �� S�  
40�� ��  S����  �  S��/  ���/���@-�$@�� 0��  S��� ����,�� 0�� �� �������@-�$0�� �� 0��  S�  ��� �� ����$�������@-�0�� 0��  S�  ��� ����(�������0��  ��0��  P� ��/���b���8@-�D0�� P��@��  T�  
�� ��k���  P�   ��8���0��4@��0�� T�����  ��8�����p@-�@�� 0��  S�p������0��  S� P��  
0��  S�  
d �吒��X0��P�� ��L0�� ��  R�  
 P��8@��  ����D���  P�p�� 0��40�� U� 0�����0�� �� ��p@�迓����j���@-� @�� ��r���  P�  
���.���  P���t �� 0��  S���  T�`@��0�40��X �� 0��a���  P�  
 �����  P�  
00��0 �� �垓�� 0��  ��0�� S�0� �  ����q���\%�Ð��j�����8@-�|P�� @�� ��  R�0�  h ��@�� @��?���  P�  
 ������  P�	  
<0��< �� ��|���  �4�� Q�0����4@�� 0��0�� ��0��0��40��8�����j���0@-��M�@�� �� P���� ������ ����b���Ѝ�0���{���s@-� @��`�� P��  T� ���� ��  
N���p ��  T� ��P��  
@�� 0��  S�@� U����|���@-�@������������ ��@������80��  P�0@-�$�M�P��  ��$�� ���@����� ��������$Ѝ�0��������ð0���@-� `��  ��  R�@� P�  � ��9���   � ��������p��P��  P�  
�� �� ��_���X0��4@�� �� T���� P��@@���� 0�� ���� ��  P�  �� 0�� �� ��  �H��� 0�� U����  ��������ώ��d2��  ���D-� @��  ���M� ��@ �㧪��D2��D"�� S�  
 ��V��  P�0��  �	  �("�� R�  
 �����  P���  �   ���	����1��@��  T�  ���P�����? �㉪��o  ���� P�㍑�� ���A �オ��  ���������������  Z�  
 ��
��?���  P�  x1���� @��ԙ�� �� ��T���  P�  
���͙��p�� ����s��� ��l�� ��)���  P�  
`��T�� �� ��"���  P�  
 ���� �����  P�  
��$��Ǚ������ę���������� ���� ������00��  S�  
�0��  U���� �� ������� ��B���  P�   ��!���  P�  
 ����0��h`��P��4@��0�� T��� ��  Q�  
� ��.���  P�  
 ������  P�  
$0��l �� ��   �` ��i���
 ����� ��Ѝ�������@����É�����ê���Ɍ��ώ������Z��X[���������@�����H���h��È��Ó���j��� 4�� ��p ���/�0�� ��  ���/����/�0�� ���/��� 0�� ��  ����0�� ��  Q�A�����"8��r ��"8��r ��r ���/�@-������?� ��0 � s�  �3��� 0��@-�" S�� B 0��   ��@� B� @��  R� ��  ����0��  \�  
" \���� 0�� 0����� 0P�@-�  ���� 0��00C�s0��	 S�� �  � ��
 �� ���p ��@�����@-黐��@������@-�,0�� ������/��? � P� � 
�� 
�� P� � ����H��@-�@������?� P�  
:C� P�   ����@��)��� *���� ��"*��@��9����I��2r��@-� ̠��, ��8 � ̌� ��Č� ��#Č�\8��\���,,�� ���������'�����蠍��@-�  ��g�� 	�� 	�������8@-� P�� @P�@�8��  ����g��@�� ��8����� �������F-�(������ @�� ���0�|p��P��  � � �� `��E0��`��p �� 0��p��Q��댐��0�� �� �� ��s ��J�����@0��`��0�� 0��0��0��	0�� �� �������� ������z ��:�����u ��7�����w ��4���a��
���� ��=���  �� ���������@-�0�� @��`��rP��� � ��#������o� �� P� `� ��`����� ��\�� �����:��#:�� S�   �����0�� ��	  �
��0��0�� 
��	��� �� �����0���� ������H�����@-� �� �� ������ �����@-� ������0��$ �� P� �  ������@-�0�� ��#������������\4�� Q��N-�p�� P��,��( �� �@�������o � ������ @��
 T� ����������
 P� ��� ���������5 � P�  ʴ��pG�@������  �P�pG@�   W��  �J��$J�� T��  
� ��pG����@�� j�������&j��	����? �)��� Y�  
 V�`
 	 V��  P�\  
8 � P��   W���\�� ��^  ڰ ����� P��  � �����P��  0�� S��  0�� S��  ���0��  S�  
p��`�� �����0�� P�  � ����� P�  
 P�    ���( � �����Q���<�� ��0���� ���
 ����� ��	������� �� �����	 ������� ����  �dB��00��  S�  
40��  S�  
 ��_���80�� P�  �� ��4 ������4�� ��< ������< ��@����� 0��40��00��@0��|  � W�z  �� ��I���  W� ���  �  �������Ѝ��N�蹗�� 0��� �@ R�k  0� S�h  � ��
��S���  P�  ���Ѝ��N�蕗����� ��,���t1��0��  S�  
 P� pU  � ��$��� i��&i��  V�O  	0�� S�;  ��p�� Q�  
 Q�  
  Q� � �0�>  
@  �0�� S�=  ����Ѝ��N�肗����� �� ��0��	��0��0�� 0����� �����	 ����� ����`��`����� �������
�� ������ 0��J���  �� �� 0�� ��`��������  �� �� ��Ѝ��N����� S�  ������� `�������� P���������� ��0@� ���������Ѝ�������H�ì�����ü������э��ߍ���A-��P��( ����D`�� �����0�� ���� @����p����0��<���� ��0����0��0��F����� ����� 0��0��0��0��0��0��0��00����H ��#� �  
L0��  S�  4 ������00��80�� ��P��8�����D ��`����A��������L�������D-�A�� �� P��P���X��`��
 �����<p��$0��+��
��4��� ��00��O���E0�� ��� 0��;��p��P�� ��0��0��0��p ��o�����@0�� �� ��0�� 0��0��	`��P������$�� ������
��
 ��m���0��  ��p �� ��1��Q��Q����0��5��T������� ��^���<0��``��
0c�0��@0�� 0�� ��s0��1���d��d ��}��� ���������N-� pQ� P��������0��� p�Q�  
1�� w�P�A�� �� ��0��X��0������ �P�$  <`����+�����4P��P�� ��0p������	0���� �� ��� `�� �����<��D0��
 ��a� ���������<0�����`c�0��`P�� ��`��@`��d��d ��B��� ��  �D`����+�� �������� ��	0�� ��� `�� �����D ��0��``���+���  ��Ѝ�����L�ä��@-����0�� ��  �������@-�� ����� @P�  
������  P�  
 ��������  P�	  
 �������  P� �  
 �� �� �����@��h0��  S�  :����  �|@��h0��0��h0������l �� p�  �3V���  ������p0��  S�0�  
t0��  ��p �� S�  
�,��B���( ��@�����0�� 0�����&���jP��\%��/��ä��$���8���@-�\@��00��  S���  ��9d��d ��3�  b� R����`0��0��`0�� S�  �  ������ 0��`0��@�����d ��@��������4���@-锍��@�����x3��x#���D-� P�� �� @�� ���M���T�X��̀�D ��`����ˀ�<��\�� ����@��X� ��l��h ��t��4��0��8��������� �����  P�  �d����B�� ���b���� ������0�� 0�� ���P����4��  S� p��  
�� �����������묢��L ��������H ��������������� ��������t�� ��	 U�0  �0��5���  ! � �  R�    �&  
02��$0��  S�  D��  �2���4��  S�4�  
2��0��  S�$�  
 �� ��������  P�  4��� p� ��  
  P�  
  ����|���j  ����y���  ���劕��%���%  �1�� ��t �� U��  ����`���`������`���0���`���\��È �  �!�� 0�� 0��H!��0��U���  �D��� ��x��m���t���~���l������a���   �h �1��  ���$��*����@������ `P�  
���8��F���5  �6���0�� ��  S�  
rc�� ��0��  b� R�  �0��`��3�/� �� 0�� S�  
 S�!  
 S����0��l0��a���xP�����  Q�  
@�� �� ��8����$���� ��g����� ��	���0���� ��  ��_����� ���������0�����Ѝ���������  �������Ü.��k-��BP��H��LP��'��_���`���e��È��ç������G��Ď�������Ì��!���L���,���2���:��� ����H ���_���, � ���8 � ����#���/�@-� @��v��� @�  ��  � 0��/ S�   ����� @� P����*���@-� @������  �� 0�� �� C�����N-�B�M�@����� `�� ��� �� p������ ��W���4��0��0��0����� ���P�� ������0��@��@�� ��	 ��p������0�� � ��  
 Y�	���K���q��	 ���� ������0��  U�P�� 0��EQ��!��1�� ����0�� ��0��0�� ��0��Bߍ�����a2��p@-��M� @��`�� ������  ����� 0�� P�  0��  S�  0��  S�  P��  U�  P0�� T�  
0�� T�0�
   �����0�� ��  � �����0�� ��   � 0�� ��ۍ�p���4�ã� 0@-��M��M� �� �� ��P�����  ��s���h0��  �� P�   ��  R�   ��  R�   ��  R�
  @��  T�  ��� ����  �������� ��   �  ��Ѝ�ۍ�0���4��@-��M� �� �� ��u���  ��N���T0��  �� P�   ��  R�   ��  R�	  @��  T�   ����  ��@��:��� ��   �  ��ۍ����4��0@-��M��M� �� �� ��P��S���  ��,���`0��  �� P�   ��  R�   ��  R�   ��  R�  @��  T�  0 ����  ��=��� ��   �  ��Ѝ�ۍ�0���4�������D-� @��  ���M��M�`�� ��P�����  �����t�� 0��p��0�� �� ������p�� �� ������  U� ��  
 ��
�� ��!�����l0��Q��P�� `������ ���� ��  �����H0�� T�o �  
< ��,0�� T� � ��� P��$ ��T0��P��%���Ѝ�ۍ�����4����à� ��  4��0@-�D�M� @��P�� @��@��@��@������ �� �������� ��0��Ġ�@����� �� �����DЍ�0��蠆 p@-��M� `��6��� @�� ������ P�� ����� � ��  
  T�0��  ��0��C1��!���� �� ������0��@�B@�Q��@�� ��P�� ��0a���C1�����ڍ�p��襆 H0��@-��M� �� r�  
0��  S�  
 ��@����� ���� 0d� ��C1��o���ڍ����4�å� �@-��M��M� p������ @�� �������  �� `����� ��$P��n��� �  ��  
  T�0��  ��0��C1��!���� �� �����0��@�B@�Q��@��$ ��P�� ��0a���C1��C���Ѝ�ڍ�����4�ã� �@-��M��M� p��`�� ��P��f���P��  �� @��i��� ��B���  �� ��?���,0��0e� �� ��(��C1����$ �� ��#���Ѝ�ڍ�����4�ã� 0@-��M��M� ��@��H���0��  �� P�� P��J���0d� �� ����C1�����Ѝ�ڍ�0���4�ã� |0��X0��0C� S��  ���ð��ü�������������������L ����  �D ����5���00��\ ��J���o��� 0��` ����� 0��  ��0��d����������/�4�å� �� T��s@-��Q���1���A�� �� 0��l ��  Q�\ ����h��P0��  �1������ ���\4��\���| �� ���,̠�������\ ��|������\��t��ޒ��  �:�� ��I��� `P�\ ��  
 �������P ��\ ������$Q��$A��\ ������` ��\ ������\ ����� ����Ē��P���� ������ �� 0��  S�  
�0�� 0��  S�  
� ��  ��  �� � 0� R�  
� �寒��0���@��� ��\��` �婒����  Q�  
��� �壒�� �� �������,���0�� �� �嚒����}����� ��&���80�� ��� ����p ��ȃ����X����Ϡ�T������Ѝ�p@��e���4��p3�È4�ü��]����<�����!��ë�������������3��	������a2��H ��3���<���\��� 4���D-��M� �� �� ���@�����  ��b���p�� 0�� P�(  0��  S�%  0��  S�"  0��  S�  P��  U�   �� ���O��� 0��/ S� `��  
`��\ ��}���\ ������ ��
�� p��\ ��`��  ��d���\0��  �
��\ �� ��^���\0�� ��P��   �  ��ۍ�����4�á��0@-��M��M� ��d �� P�� ��M���  ��&����0�� 0�� P� @�6  0��  S�2  0��  S�  0��  S�  0��  S�  
0��  S�&   ����� @`�#  �0��  ��  P�  
��� �  Q�  � ������t0����  �� �  Q�  # �㍒��` ������L0��d�� 0��  �� @��D ��P��  ��  �����40��  �� R� P�5   �$@�� ��Ѝ�ۍ�0���4��T��  ����H ��t3���������� ��@-�T0�� Q���X0��0C� S��`  ���ø�����������,��è���l��� ��d��!��� ��P  � ��T����� ��K  ���8A��B���  P�8�  0��X0��D  ���$A��`���  P�  
�妑��0��  ��墑���0��h0�� 0��������@��q���  P�  
� �嗑��0������0��X0��;��d0���0��  ��%  ���@��,���  P� ����\ �����` ��\ �����0��X0��\ ��  ���Y����� @��}�����  T�d0��  ��@�� @��
  �0�� S� ��  �  T�0� �h � ��0��X ��@��X������4�å� �� T��ä��m��Ç��Î���T�ë���<���@ ��@-�8��0��8�� S�  �( ��Q���@������ ��M���}����r���@��:���4��;���Đ��<��� 4�� ��p ���/�\1���@-� `��'���P!�� 0��0C� �� @�� S��  ����Ì��è������Ì��� @��>  �P��<����0�� ��X��� ������`����� �� p��P�� ��O������ ��L���  ����� ����  �� ��[��� ����� ���0�� ���� ��� �� P�� ��P��� P��@d�  �;��0������� ��@��  �<��t��0�� ��<��0��)���@��  �<��T��0�� ��<��0�� ���@�� �� @��4 ���� ��A����������8=��<=��X��ǐ����Å���͐��ې����� 4��s@-�h��~���  P�  
 ��
 ������P2�� ��L��u���  P�  
 ��
 ������,2��  ��$B�� ���Q�  *��א���?�� 0��b��2��B�� P�� 0��  U�0��  �1�� ����� ���\4��\���| �� ���,̠���������� �� ��������P����庐��  � ��:��%��� PP�  �� �� ������P��  � ��b����� �� �� ������ 0��0��x���XQ��PA�� ��X�埐����P�� �ᛐ��H�� 0��  S�  
<1�� 0��  S�  
  �� �� � 0� R�  
�勐��A��
 ��������児����  Q�  
���� ����� ��� ����������
 ��P������0��� �� `��@�� ��q���� ��[���0�����  ��0��~��� ������ ��`��E0��0��0�� 0��^����m � ��`�� ��;����0��O���<��1��Ѝ�p@����������X��������4��p3��8=�ü��f������!���M�������������3��<=��{������a2��H �Ê���H������t��� 4��H ��@-�D@��0����0��0�� S�  �, �����@������  �����  ����;���@������8=��X��;���Đ����Ä��D-�`�� �� @�� Q����  �� R�  
� �� V���� S������ ��PC������� P�w  
 P�  
 P����  �2�� ��
@��p��`��  ��  �O��� P�   ��
 �������1����@�� W� �����p�����:�D����� U������ �����1��  P� p�� ��  ��� �������������������!��ۏ��  � @�
���  �  Q�  # ��]���  � �� ��  �  Q�  H�巏��01��  �� R� R  ���  �� ��`�� Q�  �� �� �� ��  
�序��9  ��@��0�� �� S�����`��PE�0��
0�����  ��0���������0������@L� ��0$�0��  ��  ��@�����0��  �� R� @�5F���t0��1�� U����(� �偏�� ��  � ��8�����  ��h �协�� ��2��� @� P�  �P ��r���4��� ��D0��  ������< ��k����D�����8=��X�ß��ç��ù��ý������H ��t3�Ç���������ä�����  ���/��/� Q��/t  : P�k  � �l  
?o�/o�0B�0s�0�  ���  ��P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �
P� ���
@ 
P� ��
@ �	P� ���	@ 	P� ��	@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ �P� ���@ P� ��@ � P� ��� @  P� �� @  ���/� �  ��/�/o� b�0���/�  P�  ��  �  Q����
@-����@�� �A��/�  Q�  
� � aB Q�p  
 0�� 0`B S�o  � �q  
/o�o� @� r� �  ���  ��S�  ���?C S�  ��?C �S�  ���>C S�  ��>C �S�  ���=C S�  ��=C �S�  ���<C S�  ��<C �S�  ���;C S�  ��;C �
S�  ���:C 
S�  ��:C �	S�  ���9C 	S�  ��9C �S�  ���8C S�  ��8C �S�  ���7C S�  ��7C �S�  ���6C S�  ��6C �S�  ���5C S�  ��5C �S�  ���4C S�  ��4C �S�  ���3C S�  ��3C �S�  ���2C S�  ��2C �S�  ���1C S�  ��1C � S�  ���0C  S�  ��0C   \�  `B�/�  <�  `B�/�  �3�� ��/�/o� b�  \�3��  `B�/�  P�����+  �  Q����
@-�u���@�� �A��/� 0R� �b�0�A1�Q�A1���/� 0R� �b�0�AQ�Q�AQ���/� 0R� �b��A�Q0�A���/�  S�  R    Q�  P �  �  ��M� `-�  ����Ѝ� ���/�@-� ����������C-�@��P�� `��p��9 �������T$� ��	0��`V�p�� 0���`�������C-�@��P�� `��p��	  �������T$� ��	0��`V�p�� 0���`������  Q��O-� `���M��  �  S��  � �S����@�� P��3   R�?  �?o�  S�  c0"�C���$���S��� �������x��'x�� ��� �� ���	�%������ S�  �����I�  * S��I�����c��� ��v����� ��� ��������� X��X�� W�  �P���J�  * W��J�	��� p��  � \�B  � p�����  V�
 ��0��  
  r� 0���� ��Ѝ�����  R�  �� ��Q��� @���o�  Z�  ������d�(���$x������
 ��D����� ���
 �����	�%������ S�  �����I�  * S��I�����c��� ��1����� ��� ������8��#X��X�� X�  �P���J�  * X��J�	���p�����o�  W�  
 g�2���01�����;�����(���	��
 ��������	�� ���
 ������� �� ��� �"Ƞ�'��8�� P�  �0���K�t  :@`�	�� �� ������0��	�� @�� ��r��� ��

� (��"Ƞ� ��8�� Z�  �0��@D�[  :j����*Ƞ�"�����H�� �����������"��(�� Q�  : ����P� p��p�  W�t��
�J� p��q���  r� 0��`��0���  p� �� `��*��� pj�57��J��;�����$x���� ����������� ��� ��7���(��"�������,���8�� R�  �0���K�(  :�b���	 ���������� ��� ����"��� ��Ƞ�	�,��8�� R�  �0���I�  * R��I�0����Z������b�M��� \�  R!���0���-��� Z�0��@D����� P��K�0������ R��K�0������  S��O-�@���M� ���`�����p��P�����3   R�  �?o�  S�  c0"�S���%h������
 ��l�����H��$H�� ���
 ������	�(������
 S�  �����I�  *
 S��I����
�c���
 ��W����� p��
 �������(��"����� T�  ����pG�  * T�pG�	��� ��  � S�  �oo�  V�~  
 f�2���0��v��4������'���
�� �����5���
�� ��� �������0�� H��	�#���6����� R�  �����I�  :�b�
�� �� 0�� ���
�� P�� ���������8��#(�� 0��(�� T�  � ��PE�  :@d�	���)��#�� ���X�������������"(��,�� T�  :  � �R� �� �  Q�?  
�I� ��<  �  R�  �� ������ P���o�  Y�6  ��@e�!���%x��`���� �������� ��� ��]���	�((����� S�  �����I�  * S��I�����c��� �������� @�� ��J���

�Ƞ�,������ Z�  ����@D�  * Z�@D�	�����  � S�  R!�����  � �����	 ��Ѝ����� pi�8��Y��4g�����%x���� �������������*��� ��� ��"�������,h��H�� S�  �@���K�   :@c��� ������� `�� ����� ��� H��$8��H�� R�  �@��`F�  * R�`F�@�����@b�h����� T� ��PE�o��� R��I����W��� S��K�@������U-Boot 2010.12 (Jul 24 2014 - 15:09:03) for SMDK4412    �����������������������������������������'��/��7��>��E��L��S��Z��a��h��o��v��~�Å�Í�Õ�Ý��        �j��        ^��                                i��    �h��    lh��            4h��do_env_import   do_env_export      ������������������������������������   ����������������������������������������   set_default_env env_import  �m��n��&n��6n��@n��Ln��Vn��vn���:�ä���        �  �  �              �                          s3c_onenand_wait      *|��  2|��  :|��  B|���  J|��Z  R|��j  Z|��z  b|�Ê  j|�� �  r|��!�  z|��            �     �  ""  $I  RJ  �T  UU  U�  ��  ��  ��  ��  ��  ��  	   �   	   �	  �   �@  @  ,S E C   S 3 C 6 4 0 0 X   T e s t   B / D S y s t e m   M C U   S M D K E X Y N O S - 0 1 A n d r o i d   1 . 0 G o o g l e ,   I n c 	
 �  @   	   �   	   �	  �   �    
 �B@   �A���O�ÐO��FAT           !B c0�@�P�`�p�)�J�k���������1s2R"�R�B�r�b9��{�Z��Ӝ�����b$C4 �d�t�D�Tj�K�(�	������ō�S6r&0�v�f�V�F[�z��8�����׼��H�X�h�x@a(#8���َ��H�i�
�+��Z�J�z�jqP
3:*���˿���y�X�;���l�|�L�\",<`A�������*��h�I��~�n�^�N>2.Qp���������:�Y�x�����ʱ��-�N�o�� �0� P%@Fpg`������ڳ=���^���"�25BRwbVr�˥����n�O�,���4�$��ftGd$TDۧ������_�~��<��&�6��WfvvF4VL�m��/�ș鉊���DXeHx'h���8�(}�\�?����؛����uJTZ7jz�
��*�:.��l�Mͪ����ɍ&|ld\EL�<�,���>�]�|ߛ���ُ��n6~UNt^�.�>��    �0w,a�Q	��m��jp5�c飕d�2�����y�����җ+L�	�|�~-����d�� �jHq���A��}�����mQ���ǅӃV�l��kdz�b���e�O\�lcc=���� n;^iL�A`�rqg���<G�K���k�
����5l��B�ɻ�@����l�2u\�E���Y=ѫ�0�&: �Q�Q��aп���!#ĳV���������(�_���$���|o/LhX�a�=-f��A�vq�� Ҙ*��q���俟3Ը��x4� ��	���j-=m�ld�\c��Qkkbal�0e�N b��l{����W���ٰeP�긾�|�����bI-��|ӌeL��Xa�M�Q�:t ���0��A��Jו�=m�Ѥ����j�iC��n4F�g�и`�s-D�3_L
��|�<qP�A'�� �%�hW��o 	�f���a���^���)"�а����=�Y��.;\���l�� �������ұt9G��wҝ&���sc�;d�>jm�Zjz���	�'� 
��}D��ң�h���i]Wb��ge�q6l�knv���+ӉZz��J�go߹��ﾎC��Վ�`���~�ѡ���8R��O�g��gW����?K6�H�+�L
��J6`zA��`�U�g��n1y�iF��a��f���o%6�hR�w�G��"/&U�;��(���Z�+j�\����1�е���,��[��d�&�c윣ju
�m�	�?6�grW �J��z��+�{8���Ғ�����|!����ӆB������hn�����[&���w�owG��Z�pj��;f\��e�i�b���kaE�lx�
����T�N³9a&g��`�MGiI�wn>JjѮ�Z��f�@�;�7S���Ş��ϲG���0򽽊º�0��S���$6к���)W�T�g�#.zf��Ja�h]�+o*7������Z��-EPTGMK  0123456789abcdef    0123456789ABCDEF                             � �         	 
         # + 3 ; C S c s � � � �                                     @ @       	    ! 1 A a � � � 0@`    `   P   s   p  0  	� 
  `     	�     �  @  	�   X    	� ;  x  8  	�   h  (  	�    �  H  	�   T   � +  t  4  	�   d  $  	�    �  D  	�   \    	� S  |  <  	�   l  ,  	�    �  L  	�   R   � #  r  2  	�   b  "  	�    �  B  	�   Z    	� C  z  :  	�   j  *  	�  
  �  J  	�   V   @  3  v  6  	�   f  &  	�    �  F  	� 	  ^    	� c  ~  >  	�   n  .  	�    �  N  	� `   Q   �   q  1  	� 
  a  !  	�    �  A  	�   Y    	� ;  y  9  	�   i  )  	�  	  �  I  	�   U   +  u  5  	�   e  %  	�    �  E  	�   ]    	� S  }  =  	�   m  -  	�    �  M  	�   S   � #  s  3  	�   c  #  	�    �  C  	�   [    	� C  {  ;  	�   k  +  	�    �  K  	�   W   @  3  w  7  	�   g  '  	�    �  G  	� 	  _    	� c    ?  	�   o  /  	�    �  O  	� `   P   s   p  0  	� 
  `     	�     �  @  	�   X    	� ;  x  8  	�   h  (  	�    �  H  	�   T   � +  t  4  	�   d  $  	�    �  D  	�   \    	� S  |  <  	�   l  ,  	�    �  L  	�   R   � #  r  2  	�   b  "  	�    �  B  	�   Z    	� C  z  :  	�   j  *  	�  
  �  J  	�   V   @  3  v  6  	�   f  &  	�    �  F  	� 	  ^    	� c  ~  >  	�   n  .  	�    �  N  	� `   Q   �   q  1  	� 
  a  !  	�    �  A  	�   Y    	� ;  y  9  	�   i  )  	�  	  �  I  	�   U   +  u  5  	�   e  %  	�    �  E  	�   ]    	� S  }  =  	�   m  -  	�    �  M  	�   S   � #  s  3  	�   c  #  	�    �  C  	�   [    	� C  {  ;  	�   k  +  	�    �  K  	�   W   @  3  w  7  	�   g  '  	�    �  G  	� 	  _    	� c    ?  	�   o  /  	�    �  O  	�    A @ !  	 � @   �  a ` 1 0 � @         	  
             J���Z���a2��e���p���}��È��Ü��é���a2��              bootcmd ext3format mmc 0:3;ext3format mmc 0:4;movi read kernel 0 40008000;movi read rootfs 0 41000000 100000;bootm 40008000 41000000 vol_arm: %X
 vol_int: %X
 vol_g3d: %X
 buck1_ctrl: %X
 buck2_ctrl: %X
 buck3_ctrl: %X
 ldo14_ctrl: %X
 vol_mif: %X
 buck4_ctrl: %X
 TrustZone Enabled BSP
 BL1 version: %s
 Using half synchronizer for asynchronous bridge
 

Checking Boot Mode ...  OneNand
  NAND
  SDMMC
  EMMC4.3
  EMMC4.41
 reset... 


  select Fail. 
 Error Eint No. 
 Error Filter Width. 
 initial raw table fwbl1 u-boot parted u-boot TrustZone S/W kernel rfs bl2 
CPU: S5PC220 [Samsung SOC on SMP Platform Base on ARM CortexA9]
 APLL = %ldMHz, MPLL = %ldMHz
 This CLOCK is Not Support: %d
 

%s

 ### ERROR ### Please RESET the board ###
 Reserving %dk for malloc() at: %08lx
 Reserving %zu Bytes for Board Info at: %08lx
 Reserving %zu Bytes for Global Data at: %08lx
 DRAM:   ipaddr loadaddr bootfile Net:    bootargs machid Using machid 0x%x from environment
 [err] boot_get_ramdisk
 
Starting kernel ...

 pc : [<%08lx>]	   lr : [<%08lx>]
sp : %08lx  ip : %08lx	 fp : %08lx
 r10: %08lx  r9 : %08lx	 r8 : %08lx
 r7 : %08lx  r6 : %08lx	 r5 : %08lx  r4 : %08lx
 r3 : %08lx  r2 : %08lx	 r1 : %08lx  r0 : %08lx
 Flags: %c%c%c%c   IRQs %s  FIQs %s  Mode %s%s
 Resetting CPU ...
 fast interrupt request
 not used
 data abort
 prefetch abort
 software interrupt
 undefined instruction
 USER_26 FIQ_26 IRQ_26 SVC_26 UK4_26 UK5_26 UK6_26 UK7_26 UK8_26 UK9_26 UK10_26 UK11_26 UK12_26 UK13_26 UK14_26 UK15_26 USER_32 FIQ_32 IRQ_32 SVC_32 UK4_32 UK5_32 UK6_32 ABT_32 UK8_32 UK9_32 UK10_32 UND_32 UK12_32 UK13_32 UK14_32 SYS_32 resetting ...
 %-12s= 0x%08lX
 arch_number boot_params DRAM bank -> start -> size ethaddr (not set) %-12s= %s
 ip_addr     = %pI4
 baudrate    = %d bps
 TLB addr relocaddr reloc off irq_sp sp start  FB base   bdinfo print Board Info structure ## Starting application at 0x%08lX ...
 ## Application terminated, rc = 0x%lX
 go start application at address 'addr' addr [arg ...]
    - start application at address 'addr'
      passing 'arg' as arguments reset Perform RESET of the CPU 
## Checking Image at %08lx ...
    Legacy image found
    Bad Magic Number
    Bad Header Checksum
    Verifying Checksum ...     Bad Data CRC
 OK
 Unknown image format!
 ## Transferring control to OSE (at address %08lx) ...
 ## Transferring control to RTEMS (at address %08lx) ...
    XIP %s ...     Loading %s ...     Uncompressing %s ...  GUNZIP: uncompress, out-of-mem or overwrite error - must RESET board to recover
 Unimplemented compression type %d
 ## Transferring control to NetBSD stage-2 loader (at address %08lx) ...
 verify ## Booting kernel from Legacy Image at %08lx ...
 Unsupported Architecture 0x%x
 Wrong Image Type for %s command
 Wrong Image Format for %s command
 ERROR: can't get kernel image!
 ERROR: unknown image format type!
 Could not find kernel entry point!
 Ramdisk image is corrupt or invalid
 Trying to execute a command out of order
 initrd_start initrd_end cmdline subcommand not supported
 bdt subcommand not supported
 prep subcommand not supported
 Boot with zImage
 WARNING: legacy format multi component image overwritten
 ERROR: new format image overwritten - must RESET the board to recover
 autostart %lX filesize ERROR: booting os '%s' (%d) is not supported
 bootm boot application image from memory [addr [arg ...]]
    - boot application image stored in memory
	passing arguments 'arg ...'; when booting a Linux kernel,
	'arg' can be the address of an initrd image

Sub-commands to do part of the bootm sequence.  The sub-commands must be
issued in the order below (it's ok to not issue all sub-commands):
	start [addr [arg ...]]
	loados  - load OS image
	cmdline - OS specific command line processing/setup
	bdt     - OS specific bd_t processing
	prep    - OS specific prep before relocation or go
	go      - start OS boot default, i.e., run 'bootcmd' bootd iminfo print header information for application image addr [addr ...]
    - print header information for application image starting at
      address 'addr' in memory; this includes verification of the
      image contents (magic number, header and payload checksums) loados cmdline bdt prep OFF Data (writethrough) Cache is %s
 Instruction Cache is %s
 icache [on, off]
    - enable or disable instruction cache dcache enable or disable data cache [on, off]
    - enable or disable data (writethrough) cache List of available devices:
 %-8s %08x %c%c%c  coninfo print console devices and information echo args to console [args..]
    - echo args to console; \c suppresses newline ## No elf image at address 0x%08lx
 ## Not a 32-bit elf image at address 0x%08lx
 tftp Automatic boot of VxWorks image at address 0x%08lx ... 
 ## Ethernet MAC address not copied to NV RAM
 bootaddr eth(0,0) %s:%s  srv %s:file  e=%s  serverip h=%s  hostname tn=%s  ## Not an ELF image, assuming binary
 ## Using bootline (@ 0x%lx): %s
 ## Starting vxWorks at 0x%08lx ...
 ## vxWorks terminated
 ## Starting application at 0x%08lx ...
 ## Application terminated, rc = 0x%lx
 bootelf Boot from an ELF image in memory [-p|-s] [address]
	- load ELF image at [address] via program headers (-p)
	  or via section headers (-s) bootvx Boot vxWorks from an ELF image  [address] - load address of vxWorks ELF image. exit exit script usage : ext2format <interface> <dev[:part]>
 
** Invalid boot device **
 
** Invalid boot device, use 'dev[:part]' **
 ** Partition Number shuld be 1 ~ 4 **
 Start format MMC%d partition%d ....
 Format failure!!!
 FileSystem Type Value is not invalidate=%d 
 ** No boot file defined **
 ** Bad partition %d **
 U-Boot ** Invalid partition type "%.32s" (expect "U-Boot")
 Loading file "%s" from %s device %d:%d (%.32s)
 Loading file "%s" from %s device %d
 ** Bad partition - %s %d:%d **
 ** Bad ext2 partition or disk - %s %d:%d **
 ** File not found %s
 %d bytes read
 %X 
** Block device %s %d not supported
 
** Invalid boot device, use `dev[:part]' **
 / ** Error ext2fs_ls() **
 ext2ls list files in a directory (default /) <interface> <dev[:part]> [directory]
    - list files from 'dev' on 'interface' in a 'directory' ext2load load binary file from a Ext2 filesystem <interface> <dev[:part]> [addr] [filename] [bytes]
    - load binary file 'filename' from 'dev' on 'interface'
      to address 'addr' from ext2 filesystem ext2format ext2format - disk format by ext2
 <interface(only support mmc)> <dev:partition num>
    - format by ext2 on 'interface'
 ext3format ext3format - disk format by ext3
 <interface(only support mmc)> <dev:partition num>
    - format by ext3 on 'interface'
 [Partition table on  OneNAND MoviNAND ptn %d name='%s'  start=0x%X  start=N/A  len=0x%X(~%dKB)  len=N/A  (Yaffs)
 (use hard-coded info. (cmd: movi))
 fbparts Fastboot: Adding partitions from environment
 Error:FASTBOOT size of parition is 0
 Error:FASTBOOT offset of parition is not given
 Error:FASTBOOT no partition name for '%s'
 Error:FASTBOOT no closing %c found in partition name
 yaffs swecc hwecc Error:FASTBOOT partition name is too long
 Error:FASTBOOT no name
 Error:Fastboot: Abort adding partitions
 Fastboot: employ default partition information
 No partition informations! Adding: %s, offset 0x%8.8x, size 0x%8.8x, flags 0x%8.8x
 Error: Image size is larger than partition size!
 flashing '%s'
 write mmc %d Compressed ext4 image
 *** erase start block 0x%x ***
 *** erase block length 0x%x ***
 erase user mmc %s %s %s %s %s
 *** erase block length too small ***
 zero emmc open 0 tzsw rootfs emmc close 0 userdata fat Error: No MBR is found at SD/MMC.
 Hint: use fdisk command to make partitions.
 flash undefined image name !
 Fastboot inactivity timeout %ld seconds
 Fastboot ended by user
 Fastboot error 
 Fastboot disconnect detected
 Fastboot inactivity detected
 No variables set ERROR OKAY 
downloading of %d bytes finished
 Warning empty download buffer
 Ignoring
 FAIL reboot -bootloader getvar: 0.4 product serialno downloadsize erase: FAILpartition does not exist erasing(formatting) '%s'
 erasing '%s'
 ext3format mmc 0:3 ext3format mmc 0:4 fatformat mmc 0:1 FAILfailed to erase partition partition '%s' erased
 download: Starting download of %d bytes
 FAILdata invalid size FAILdata too large DATA%08x Kernel size: %08x
 Ramdisk size: %08x
 Booting kernel..
 setenv Booting raw image..
 ERROR : bootting failed
 You should reset the board
 FAILinvalid boot image flash: FAILno image downloaded FAILimage too large for partition flashing '%s' failed
 kernel+ramdisk FAILfailed to flash partition partition '%s' flashed
 Unknown Error savenv '%s' failed : %s
 FAIL%s partition '%s' saveenv-ed
 oem INFOunknown OEM command fastboot fastboot- use USB Fastboot protocol
 [inactive timeout]
    - Run as a fastboot usb device.
    - The optional inactive timeout is the decimal seconds before
    - the normal console resumes
 usage : fatformat <interface> <dev[:part]>
 
 ** Invalid boot device **
 
 ** Invald boot device, use 'dev[:part]' **
 ** Partition Number should be 1 ~ 4 **
 Start format MMC&d partition&d ...
 usage: fatinfo <interface> <dev[:part]>
 -----Partition %d-----
 
** Unable to use %s %d:%d for fatinfo **
 ------------------------
 usage: fatls <interface> <dev[:part]> [directory]
 
** Unable to use %s %d:%d for fatls **
 No Fat FS detected
 usage: fatload <interface> <dev[:part]> <addr> <filename> [bytes]
 MMC init is failed.
 
** Unable to use %s %d:%d for fatload **
 
** Unable to read "%s" from %s %d:%d **
 
%ld bytes read
 fatload fatload - load binary file from a dos filesystem
 <interface> <dev[:part]>  <addr> <filename> [bytes]
    - load binary file 'filename' from 'dev' on 'interface'
      to address 'addr' from dos filesystem fatls fatinfo fatinfo - print information about filesystem <interface> <dev[:part]>
    - print information about filesystem from 'dev' on 'interface'
 fatformat fatformat - disk format by FAT32
 <interface(only support mmc)> <dev:partition num>
	- format by FAT32 on 'interface'
 help print command description/usage 
	- print brief description of all commands
help command ...
	- print detailed usage of 'command' ? alias for 'help' Unknown operator '%s'
 Invalid data width specifier
 -lt < -gt -eq == -ne != <> -ge >= -le <= itest return true/false on integer compare [.b, .w, .l, .s] [*]value1 <op> [*]value2 ## Total Size      = 0x%08x = %d Bytes
 ## Switch baudrate to %d bps and press ENTER ...
 loady ## Ready for binary (ymodem) download to 0x%08lX at %d bps...
 ## Ready for binary (kermit) download to 0x%08lX at %d bps...
 ## Binary (kermit) download aborted
 ## Start Addr      = 0x%08lX
 ## Switch baudrate to %d bps and press ESC ...
 
## First Load Addr = 0x%08lX
## Last  Load Addr = 0x%08lX
## Total Size      = 0x%08lX = %ld Bytes
 loads_echo ## Ready for S-Record download ...
 ## S-Record download aborted
 loads load S-Record file over serial line [ off ]
    - load S-Record file over serial line with offset 'off' loadb load binary file over serial line (kermit mode) [ off ] [ baud ]
    - load binary file over serial line with offset 'off' and baudrate 'baud' load binary file over serial line (ymodem mode) CRC32 for %08lx ... %08lx ==> %08lx
 Base Address: 0x%08lx
 Tested %d iteration(s) with %lu errors.
 Pattern %08lX  Writing...%12s Reading... 
Mem error @ 0x%08X: found %08lX, expected %08lX
 Zero length ???
 word at 0x%08lx (0x%08lx) != word at 0x%08lx (0x%08lx)
 halfword at 0x%08lx (0x%04x) != halfword at 0x%08lx (0x%04x)
 byte at 0x%08lx (0x%02x) != byte at 0x%08lx (0x%02x)
 byte halfword Total of %ld %s%s were the same
 %08lx:  %04x  %02x  ?  memory display [.b, .w, .l] address [# of objects] mm memory modify (auto-incrementing address) [.b, .w, .l] address nm memory modify (constant address) mw memory write (fill) [.b, .w, .l] address value [count] cp memory copy [.b, .w, .l] source target count cmp memory compare [.b, .w, .l] addr1 addr2 count crc32 checksum calculation address count [addr]
    - compute CRC32 checksum [save at addr] base print or set address offset 
    - print address offset for memory commands
base off
    - set address offset for memory commands to 'off' loop infinite loop on address range [.b, .w, .l] address number_of_objects mtest simple RAM read/write test [start [end [pattern [iterations]]]] sleep delay execution for some time N
    - delay execution for N seconds (N is _decimal_ !!!) Card NOT detected or Init Failed!!
 Device: %s
 Manufacturer ID: %x
 OEM: %x
 Name: %c%c%c%c%c 
 Tran Speed: %d
 Rd Block Len: %d
 %s version %d.%d
 No Yes High Capacity: %s
 Size: %dMB (block: %d)
 4-bit 8-bit 4-bit DDR 1-bit 8-bit DDR Bus Width: %s
 Boot Partition Size: %d KB
 rescan Usage:
%s
 list Default erase user partition
 Block count is Too BIG!!
 Erase all from %d block
 MMC erase Success.!!
 MMC erase Failed.!!
 read 
MMC read: dev # %d, block # %d, count %d ...  %d blocks read: %s
 OK 
MMC write: dev # %d, block # %d, count %d ...  %d blocks written: %s
 eMMC boot partition Size is %d MB.!!
 eMMC RPMB partition Size is %d MB.!!
 eMMC boot partition Size change Failed.!!
 open eMMC OPEN Success.!!
 			!!!Notice!!!
 !You must close eMMC boot Partition after all image writing!
 !eMMC boot partition has continuity at image writing time.!
 !So, Do not close boot partition, Before, all images is written.!
 eMMC OPEN Failed.!!
 close eMMC CLOSE Success.!!
 eMMC CLOSE Failed.!!
 mmcinfo mmcinfo <dev num>-- display MMC info emmc Open/Close eMMC boot Partition emmc open <device num> 
emmc close <device num> 
emmc partition <device num> <boot partiton size MB> <RPMB partition size MB>
 MMC sub system read <device num> addr blk# cnt
mmc write <device num> addr blk# cnt
mmc rescan <device num>
mmc erase <boot | user> <device num> <start block> <block count>
mmc list - lists available devices mmc/sd device is NOT founded.
 partion #    size(MB)     block start #    block count    partition_Id 
    1        %6d         %8d        %8d          0x%.2X 
    2        %6d         %8d        %8d          0x%.2X 
    3        %6d         %8d        %8d          0x%.2X 
    4        %6d         %8d        %8d          0x%.2X 
 fdisk is completed
 -c -p Usage:
fdisk <-p> <device_num>
 fdisk <-c> <device_num> [<sys. part size(MB)> <user data part size> <cache part size>]
 fdisk fdisk	- fdisk for sd/mmc.
 -c <device_num>	- create partition.
fdisk -p <device_num> [<sys. part size(MB)> <user data part size> <cache part size>]	- print partition information
 mmcinfo %d reading writing %s FWBL1 ..device %d Start %ld, Count %ld  mmc %s %d 0x%lx 0x%lx 0x%lx %s BL2 ..device %d Start %ld, Count %ld  %s bootloader..device %d Start %ld, Count %ld  %s kernel..device %d Start %ld, Count %ld  %s RFS..device %d Count %ld, Start %ld  %s %d TrustZone S/W.. Start %ld, Count %ld  movi movi	- sd/mmc r/w sub system for SMDK board init - Initialize moviNAND and show card info
movi read zero {fwbl1 | u-boot} {device_number} {addr} - Read data from sd/mmc
movi write zero {fwbl1 | u-boot} {device_number} {addr} - Read data from sd/mmc
movi read {u-boot | kernel} {device_number} {addr} - Read data from sd/mmc
movi write {fwbl1 | u-boot | kernel} {device_number} {addr} - Write data to sd/mmc
movi read rootfs {device_number} {addr} [bytes(hex)] - Read rootfs data from sd/mmc by size
movi write rootfs {device_number} {addr} [bytes(hex)] - Write rootfs data to sd/mmc by size
movi read {sector#} {device_number} {bytes(hex)} {addr} - instead of this, you can use "mmc read"
movi write {sector#} {device_number} {bytes(hex)} {addr} - instead of this, you can use "mmc write"
 nor onenand invalid partition number %d for device %s%d (%s)
 mtddevnum mtddevname %ug %um %uk %u %s%d,%d cannot add second partition at offset 0
 incorrect device type in %s
 incorrect device number in %s
 no partition number specified
 unexpected trailing character '%c'
 no such device %s%d
 no such partition
 %s%d Device %s not found!
 %s: offset %08x beyond flash size %08x
 %s%d: partition (%s) size too big
 %s: partitioning exceeds flash size
 %s%d: partition (%s) start offsetalignment incorrect
 %s%d: partition (%s) size alignment incorrect
 %s%d: partition (%s) start offset alignment incorrect
 partition size too small (%lx)
 no closing ) found in partition name
 empty partition name
 no partitions allowed after a fill-up partition
 unexpected character '%c' at the end of partition
 out of memory
 0x%08lx@0x%08lx no partitions for device %s%d (%s)
 unexpected character '%c' at the end of device
 invalid mtd device '%.*s'
 mtdids mtdparts mtdids not defined, no default present
 mtdids too long (> %d)
 mtdparts variable not set, see 'help mtdparts'
 mtdparts too long (> %d)
 mtdids: incorrect <dev-num>
 mtdids: no <mtd-id> identifier
 device id %s%d redefined, please correct mtdids variable
 could not initialise device list
 mtdparts= mtdparts variable doesn't start with 'mtdparts='
 device %s%d redefined, please correct mtdparts variable
 mtdparts_init: no valid partitions
 no partition id specified
 partition changed to %s%d,%d
 default delall 
device %s%d <%s>, # parts = %d
  #: name		size		offset		mask_flags
 %2d: %-20s0x%08x	0x%08x	%d
 no partitions defined
 
active partition: %s%d,%d - (%s) 0x%08x @ 0x%08x
 could not get current partition info

 
defaults:
 mtdids  : %s
 none mtdparts:  add no such device %s defined in mtdids variable
 too long partition description
 %s:%s(%s)%s generated mtdparts too long, reseting to null
 del current partition deleted, resetting current to 0
 partition %s not found
 chpart change active partition part-id
    - change active partition (e.g. part-id = nand0,1) define flash/nand partitions 
    - list partition table
mtdparts delall
    - delete all partitions
mtdparts del part-id
    - delete partition (e.g. part-id = nand0,1)
mtdparts add <mtd-dev> <size>[@<offset>] [<name>] [ro]
    - add partition
mtdparts default
    - reset partition table to defaults

-----

this command uses three environment variables:

'partition' - keeps current partition identifier

partition  := <part-id>
<part-id>  := <dev-id>,part_num

'mtdids' - linux kernel mtd device id <-> u-boot device id mapping

mtdids=<idmap>[,<idmap>,...]

<idmap>    := <dev-id>=<mtd-id>
<dev-id>   := 'nand'|'nor'|'onenand'<dev-num>
<dev-num>  := mtd device number, 0...
<mtd-id>   := unique device tag used by linux kernel to find mtd device (mtd->name)

'mtdparts' - partition list

mtdparts=mtdparts=<mtd-def>[;<mtd-def>...]

<mtd-def>  := <mtd-id>:<part-def>[,<part-def>...]
<mtd-id>   := unique device tag used by linux kernel to find mtd device (mtd->name)
<part-def> := <size>[@<offset>][<name>][<ro-flag>]
<size>     := standard linux memsize OR '-' to denote all remaining space
<offset>   := partition start offset within the device
<name>     := '(' NAME ')'
<ro-flag>  := when set to 'ro' makes partition read-only (not used, passed to kernel) ping failed; host %s is not alive
 host %s is alive
 gatewayip netmask rootpath dnsip domain yes Automatic boot of image at addr 0x%08lX ...
 bootp boot image via network using BOOTP/TFTP protocol [loadAddress] [[hostIPaddr:]bootfilename] tftpboot boot image via network using TFTP protocol nfs boot image via network using NFS protocol ping send ICMP ECHO_REQUEST to network host pingAddress Not implemented yet
 ## Warning: defaulting to text format
 ## Warning: Input data exceeds %d bytes - truncated
 ## Info: input data size = %zd = 0x%zX
 ## Error: bad CRC, import failed
 ERROR: Environment import failed: errno = %d

at %s:%d/%s()
 cmd_nvedit.c ## %s: only one of "-b", "-c" or "-t" allowed
 -f ## Resetting to default environment
 env_buf too small [%d]
 Saving Environment to %s...
 %s=%s
 
Environment size: %d/%ld bytes
 ## Error: "%s" not defined
 ## Error: illegal character '=' in variable name "%s"
 stdin stdout stderr Can't delete "%s"
 baudrate ## Can't malloc %d bytes
 ## Error inserting "%s" variable, errno=%d
 ## Baudrate %d bps not supported
 ERROR: Cannot export environment: errno = %d

at %s:%d/%s()
 %zX edit:  saveenv save environment variables to persistent storage environment handling commands default -f - reset default environment
env edit name - edit environment variable
env export [-t | -b | -c] addr [size] - export environmnt
env import [-d] [-t | -b | -c] addr [size] - import environmnt
env print [name ...] - print environment
env run var [...] - run commands in an environment variable
env save - save environment
env set [-f] name [arg ...]
 editenv edit environment variable name
    - edit environment variable 'name' printenv print environment variables 
    - print values of all environment variables
printenv name ...
    - print value of environment variable 'name' set environment variables name value ...
    - set environment variable 'name' to 'value ...'
setenv name
    - delete environment variable 'name' run run commands in an environment variable var [...]
    - run the commands in the environment variable(s) 'var' delete edit export import print save reginfo print register information Bad magic number
 Bad header crc
 Bad data crc
 Bad image type
 Empty Script
 Wrong image format for "source" command
 ## Executing script at %08lx
 source run script from memory [addr]
	- run script starting at addr
	- A valid image header must be present -o -a -z -n minimal test like /bin/sh [args..] false do nothing, unsuccessfully true do nothing, successfully Audio See Interface Communication Human Interface Printer Mass Storage Hub CDC Data Vendor specific Out In      - Endpoint %d %s  Control Isochronous Interrupt  MaxPacket %d  Interval %dms Human Interface, Subclass:  None Boot  Keyboard Mouse reserved Mass Storage,  RBC  SFF-8020i (ATAPI) QIC-157 (Tape) UFI SFF-8070 Transp. SCSI Command/Bulk Command/Bulk/Int Bulk only  %s +- %d  480 Mb/s 12 Mb/s 1.5 Mb/s  %s (%s, %dmA)
  %s  %s %s %s
 %d: %s,  USB Revision %x.%x
  - %s %s %s
  - Class:   - Class: (from Interface) %s
  - PacketSize: %d  Configurations: %d
  - Vendor: 0x%04x  Product 0x%04x Version %d.%d
 String: "%s"      Interface: %d
      - Alternate Setting %d, Endpoints: %d
      - Class       -     Configuration: %d
 Bus Powered  Self Powered  Remote Wakeup     - Interfaces: %d %s%s%dmA
 (Re)start USB...
 stop stopping USB..
 USB is stopped. Please issue 'usb start' first.
 tree 
Device Tree:
 inf config for device %d
 *** NO Device avaiable ***
 usb USB sub-system reset - reset (rescan) USB controller
usb  tree  - show USB device tree
usb  info [dev] - show available USB devices Now, Waiting for DNW to transmit data
 dnw dnw     - initialize USB device and ready to receive for Windows server (specific)
 [download address]
 print monitor version ## Copying part %d from legacy image at %08lx ...
 Must specify load address for %s command with compressed image
 Bad Image Part
 Invalid image type for imxtract
    Loading part %d ...     Uncompressing part %d ...  GUNZIP ERROR - image not loaded
 %8lx fileaddr imxtract extract a part of a multi-image addr part [dest]
    - extract <part> from legacy image at <addr> and copy to <dest> %s - %s

 Usage:
%s  - No additional help available.
 %-*s- %s
 Unknown command '%s' - try 'help' without arguments for list of all known commands

 In:     No input devices available!
 Out:    No output devices available!
 Err:    No error devices available!
 Invalid Version Info! 0x%2x
 Invalid File Header Size! 0x%8x
 Invalid Chunk Header Size! 0x%8x
 Invalid Block Size! 0x%8x
 Invalid Volume Size! Image is bigger than partition size!
 partion size %lld , image size %d 
 mmc write 0 0x%x 0x%x 0x%x *** fill_chunk ***
 *** unknown chunk type ***
 *** Warning - using default environment

 *** Error - default environment is too large

 Cannot export environment Unknown boot device
 SMDK bootable device *** Warning - %s, using default environment

 Using default environment

 env_common.c !bad CRC ERROR: Cannot import environment: errno = %d

at %s:%d/%s()
 !import failed syntax error
 
 ** Abort
 HUSH_VERSION 0.01 ERROR : memory not allocated
 SMDK4412 #  %s: readonly variable ERROR: There is a global environment variable with the same name.
 IFS  	
 \$'" ;&|# *?[\ ;$&| exit not allowed from main input shell.
 <INTERRUPT>
 Unknown command '%s' - try 'help' or use 'run' command
 Unknown command '%s' - try 'help'
 'bootd' recursion detected
 showvar print local hushshell variables 
    - print values of all hushshell variables
showvar name ...
    - print value of hushshell variable 'name' then elif else fi for while until do done Unknown OS Unknown Architecture Unknown Image Unknown Compression bootm_low %d Bytes =  %sImage Name:   %.*s
 %sImage Type:    %s %s %s (%s)
 %sData Size:     %sLoad Address: %08x
 %sEntry Point:  %08x
 %sContents:
 %s   Image %d:  %s    Offset = 0x%08lx
 initrd_high ramdisk - allocation error
    Loading Ramdisk to %08lx, end %08lx ...  bootm_size ## Loading init Ramdisk from Legacy Image at %08lx ...
 No Linux %s Ramdisk Image
 Wrong Ramdisk Image Format
 ## Loading init Ramdisk from multi component Legacy Image at %08lx ...
 uncompressed bzip2 bzip2 compressed gzip gzip compressed lzma lzma compressed lzo lzo compressed Invalid Image Filesystem Image firmware Firmware Kernel Image multi Multi-File Image RAMDisk Image Script standalone Standalone Program flat_dt Flat Device Tree kwbimage Kirkwood Boot Image imximage Freescale i.MX Boot Image Invalid ARCH alpha Alpha arm ARM Intel x86 ia64 IA64 m68k M68K microblaze MicroBlaze mips MIPS mips64 MIPS 64 Bit nios2 NIOS II powerpc PowerPC ppc s390 IBM S390 SuperH sparc SPARC sparc64 SPARC 64 Bit blackfin Blackfin avr32 AVR32 Invalid OS linux Linux netbsd NetBSD Enea OSE rtems RTEMS qnx QNX vxworks VxWorks ** Too many args (max. %d) **
 ## Command too long!
 %.*s %*s 
 bootdelay Hit any key to stop autoboot: %2d  %2d  serial ERROR: USB_MAX_HUB (%d) reached
 ERROR, too many USB Devices, max=%d
  ERROR: NOT USB_CONFIG_DESC %x
 selecting invalid interface %d unable to get descriptor, error %lX
 config descriptor too short (expected %i, got %i)
 cannot reset port %i!?
 usb_new_device:cannot locate device's port.
 
     Couldn't reset port %i
 
      USB device not accepting new address (error=%lX)
 unable to get device descriptor (error=%d)
 USB device descriptor short read (expected %i, got %i)
 failed to set default configuration len %d, status %lX
 No USB Device found
 %d USB Device(s) found
 USB:    scanning bus for devices...  Error, couldn't init Lowlevel part
 Unknown error Cksum xyzModem - %s mode, %d(SOH)/%d(STX)/%d(CAN) packets, %d retries
 Block sequence error CRC/checksum error Invalid framing Cancelled End of file Timed out Sorry, zModem not available yet Can't access file 
Partition Map for  IDE SATA ATAPI USB DOC UNKNOWN  device %d  --   Partition Type: %s

 DOS ## Unknown partition table
 (%d:%d) Vendor: %s Prod.: %s Rev: %s
 Model: %s Firm: %s Ser#: %s
 Vendor: %s Rev: %s Prod: %s
 device type DOC
 device type unknown
 Unhandled device type: %i
             Type:  Removable  Hard Disk CD ROM Optical Device Tape # %02X #             Capacity: %ld.%ld MB = %ld.%ld GB (%ld x %ld)
             Capacity: not available
 ** Can't read partition table on %d:%d **
 bad MBR sector signature 0x%02x%02x
 hd%c%d sd%c%d usbd%c%d docd%c%d xx%c%d FAT FAT32  Extd %5d		%10d	%10d	%2x%s
     1		         0	%10ld	%2x
 Partition     Start Sector     Num Sectors     Type
 START: %d BLOCK: %d
 high_capacity: %d
 Capacity: %d
 
Erase
 
			*** NOTICE ***
 *** High Capacity(higher than 2GB) MMC's erase minimum size is 512KB ***
 
 %d KB erase Done
 
 %d.%d MB erase Done
 
 %d.%d GB erase Done
 
 %d B erase Done
 %s: %d MMC Device %d not found
 # Tx: Inverter delay / Rx: Inverter delay
 ## Tx: Basic delay / Rx: Inverter delay
 ## Tx: Inverter delay / Rx: Basic delay
 ### Tx: Basic delay / Rx: Basic delay
 # Tx: Disable / Rx: Basic delay
 ## Tx: Disable / Rx: Inverter delay
 ### Tx: Basic delay / Rx: Disable
 ### Tx: Inverter delay / Rx: Disable
 S5P_MSHC 
count: %d
 CMD reset
 CMD Reset is NEVER released
 DATA reset
 DATA Reset is NEVER released
 

mmc write failed ERROR: %d
 data.dest: 0x%08x
 data.blocks: %d
 data.blocksize: %d
 MMC_DATA_WRITE
 mmc write failed
 mmc read failed ERROR: %d
 MMC_DATA_READ
 mmc read failed
 Could not allocate buffer for MMC read!
 unrecognised CSD structure version %d
 could not allocate a buffer to receive the ext_csd.
 unable to read EXT_CSD on a possible high capacity card. Card will be ignored.
 unable to read EXT_CSD, performance might suffer.
 unrecognised EXT_CSD structure version %d
 card is mmc v4 but doesn't support any high-speed modes.
 NAME: %s
 Man %06x Snr %08x %c%c%c%c%c MMC Device %d: %d MB
 Internal clock never stabilised.
 Controller never released inhibit bit(s).
 FAIL: waiting for status update.
 error: %08x cmd %d
 FAIL: card is still busy
 error during transfer: 0x%08x
 SDHCI_INT_DMA_END
 S3C_HSMMC%d mmc: Reset 0x%x never completed.
 Clock %s has been failed.
  Changing clock has been failed.
  Reset FIFO never completed.
 Count: %d
 Controller never released 				data0 before reset ciu.
 Reset CTRL never completed.
 Reset DMA never completed.
 Controller never released data busy!!
 there are pending interrupts 0x%08x
 [ERROR] CMD busy. current cmd %d. last cmd reg 0x%x
 [ERROR] response error : %08x cmd %d
 unexpected condition 0x%x
 [ERROR] response timeout error : %08x cmd %d
 S5P_MSHC%d REVISION: %d.%d
 U-Boot BUG at %s:%d!
 mtdcore.c Removing MTD device #%d (%s) with use count %d
 block %d is write-protected!
 %s: ECC error = 0x%04x
 %s: controller error = 0x%04x
 %s: it's locked error = 0x%04x
 s3c_onenand_writew: Illegal access at reg 0x%x, value 0x%x
 s3c_onenand_readw:  Illegal access at reg 0x%x, value 0x%x
 smc911x: Invalid chip endian 0x%08lx
 %s-%hu smc911x smc911x: Unknown chip ID %04lx
 TX_STS_LOC  TX_STS_LATE_COLL  TX_STS_MANY_COLL  TX_STS_MANY_DEFER  TX_STS_UNDERRUN smc911x: failed to send packet: %s%s%s%s%s
 smc911x: dropped bad packet. Status: 0x%08x
 %s: timeout in RX
 smc911x: timeout waiting for PM restore
 smc911x: reset timeout
 smc911x: detected %s controller
 smc911x: phy initialized
 smc911x: autonegotiation timed out
 smc911x: MAC %pM
 LAN9115 LAN9116 LAN9117 LAN9118 LAN9211 LAN9215 LAN9216 LAN9217 LAN9218 LAN9220 LAN9221 Checksum is being calculated. 
Checksum O.K.
 
Checksum Value => MEM:%x DNW:%x
 Checksum failed.

 [s3c_usb_print_pkt: %x, ---------ERROR: DMA Address is not aligned by 8---------
 Download Done!! Download Address: 0x%x, Download Filesize:0x%x
 **** Error:Neither High_Speed nor Full_Speed
 OTG cable Connected!
 Insert a OTG cable into the connector!
 Error : Current Mode is Host
 Samsung S.LSI smdk dieid# SLSI0123 Android Fastboot ERROR: index > length
 ERROR: sohci_submit_job: EPIPE
 ERROR: ep_add_ed: pending delete
 ERROR: sohci_submit_job: ENOMEM
 ERROR: need %d TDs, only have %d
 ERROR: sohci_submit_job: EINVAL
 ** Can't read from device %d **
 ** MBR is broken **
 ** Partition%d is not ext2 file-system %d **
 Partition%d: Start Address(0x%x), Size(0x%x)
 Can't make img buffer~~!!
 Can't make img2 buffer~~!!
 Can't make reserve_img buffer~~!!
 Can't make img3 buffer~~!!
 Can't make img4 buffer~~!!
 Can't make zero buffer~~!!
 Can't make img5 buffer~~!!
 Can't make rootdata buffer~~!!
 Can't make inodedata buffer~~!!
 Can't make inodedata2 buffer~~!!
 Start ext2format...
 Wirte %d/%dblock-group
 Reserved blocks for jounaling : %d
 Start write addr : 0x%x
 Can't write Superblock(%d)~~~!!!
 Can't write Descriptor Table(%d)~~~!!!
 Can't write reserve(%d)~~~!!!
 Can't write inode bitmap(%d)~~~!!!
 Erase inode table(%d) - 0x%x Can't erase inode table(%d)~~~!!!
 Can't write rootdata~~~!!!
 Can't write root+1~~~!!!
 Can't write 7th inode~~~!!!
 Can't write 8th inode~~~!!!
 Can't  inodeval~~~!!!
 d_indirect_point:0x%x
 Can't write inode table(%d)~~~!!!
 Failed to mount ext2 filesystem...
 ** ext2fs read block (indir 1) malloc failed. **
 ** ext2fs read block (indir 1) failed. **
 ** ext2fs read block (indir 2 1) malloc failed. **
 ** ext2fs read block (indir 2 1) failed. **
 ** ext2fs read block (indir 2 2) malloc failed. **
 ** ext2fs read block (indir 2 2) failed. **
 ** ext2fs doesn't support tripple indirect blocks. **
 <DIR>  <SYM>         < ? >  %10d %s
 ** Can not find directory. **
  ** ext2fs_devread() read outside partition sector %d
 ** Invalid Block Device Descriptor (NULL)
  ** ext2fs_devread() read error **
  ** ext2fs_devread() read error - block
  ** ext2fs_devread() read error - last part
 FAT32    FAT12    FAT16    No current device
 Interface:   SD/MMC Unknown 
  Device %d:  
No valid FAT fs found
 Partition %d: Filesystem: %s "%s"
 Invalid FAT entry
             %s%c
  %8ld   %s%c
 
%d file(s), %d dir(s)

 Error reading cluster
 reading %s
 ** Partition %d not valid on device %d **
 Can't erase reserved sector~~~!!!
 SAMSUNG size checking ...
 Can't format less than 32Mb partition!!
 Under 64M
 Under 128M
 Under 256M
 Under 8G
 Under 16G
 16G~
 write FAT info: %d
 Fat size : 0x%x
 NO NAME  Can't write PBR~~~!!!
 Can't make img buffer~~(reserved)!!
 Can't write reserved region~~~!!!
 Can't make dummy buffer~~!!
 Erase FAT region Can't erase FAT region~~!!!
 Can't write FAT~~~!!!
 Partition%d format complete.
 Can't load file without a filesystem!
 %s/%s Can't list files without a filesystem!
 %llu Bytes%s %lu  %ciB%s  %0*x     %s
 1.2.3 Error: inflateInit2() returned %d
 Error: inflate() returned %d
 Error: Bad gzipped data
 Error: gunzip out of data in header
 himport_r: can't insert "%s=%s" into hash table
 ERROR: Failed to allocate 0x%lx bytes below 0x%lx.
 %ld .%03ld <NULL> (null) invalid distance too far back invalid distance code invalid literal/length code incorrect header check unknown compression method invalid window size unknown header flags set header crc mismatch invalid block type invalid stored block lengths too many length or distance symbols invalid code lengths set invalid bit length repeat invalid literal/lengths set invalid distances set incorrect data check incorrect length check need dictionary stream end file error stream error data error insufficient memory buffer error incompatible version *** WARNING: %s is too long (%d - max: %d) - truncated
 Host Name Root Path NIS Domain Name autoload NFS BOOTP broadcast %d
 
Retry count exceeded; starting again
 unknown ethact ethrotate %pM eth%daddr Board Net Initialization Failed
 CPU Net Initialization Failed
 Net Initialization Skipped
 ethprime  [PRIME] 
Warning: eth device name has a space!
 
Warning: %s MAC addresses don't match:
 Address in SROM is         %pM
 Address in environment is  %pM
 ethmacskip eth%dmacskip %d.%d.%d.%d bad length %d < %d
 len bad %d < %d
 checksum bad
  ICMP Host Redirect to %pI4  ## Warning: gatewayip needed but not set
 netretry once 
ARP Retry count exceeded; starting again
 nvlan *** ERROR: ping address not given
 *** ERROR: `serverip' not set
 *** ERROR: `ipaddr' not set
 *** ERROR: No ethernet found.
 *** ERROR: `ethaddr' not set
 *** ERROR: `eth%daddr' not set
 Using %s device
 
Abort
 Bytes transferred = %ld (%lx hex)
 /nfsroot/%02lX%02lX%02lX%02lX.img *** Warning: no boot file name; using '%s'
 File transfer via NFS from server %pI4; our IP address is %pI4 ; sending through gateway %pI4 
Filename '%s/%s'.  Size is 0x%x Bytes =  
Load address: 0x%lx
Loading: * *** ERROR: Cannot mount
 *** ERROR: Cannot umount
 
done
 *** ERROR: File lookup fail
 *** ERROR: Symlink fail
 T  octet blksize%c%d%c File too large File has bad magic tftpblocksize tftptimeout TFTP timeout (%ld ms) too low, set minimum = 1000 ms
 TFTP from server %pI4; our IP address is %pI4 Filename '%s'. Load address: 0x%lx
 blksize 
	 %lu MB received
	  
TFTP error: First block is not block 1 (%ld)
Starting again

 
TFTP error: '%s' (%d)
 Not retrying...
 ���   
   	                                             ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������     0 @ P ` p � � � � � � � �   0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p�������� 		 	0	@	P	`	p	�	�	�	�	�	�	�	�	 

 
0
@
P
`
p
�
�
�
�
�
�
�
�
  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 @@ @0@@@P@`@p@�@�@�@�@�@�@�@�@ AA A0A@APA`ApA�A�A�A�A�A�A�A�A BB B0B@BPB`BpB�B�B�B�B�B�B�B�B CC C0C@CPC`CpC�C�C�C�C�C�C�C�C DD D0D@DPD`DpD�D�D�D�D�D�D�D�D EE E0E@EPE`EpE�E�E�E�E�E�E�E�E FF F0F@FPF`FpF�F�F�F�F�F�F�F�F GG G0G@GPG`GpG�G�G�G�G�G�G�G�G HH H0H@HPH`HpH�H�H�H�H�H�H�H�H II I0I@IPI`IpI�I�I�I�I�I�I�I�I JJ J0J@JPJ`JpJ�J�J�J�J�J�J�J�J KK K0K@KPK`KpK�K�K�K�K�K�K�K�K LL L0L@LPL`LpL�L�L�L�L�L�L�L�L MM M0M@MPM`MpM�M�M�M�M�M�M�M�M NN N0N@NPN`NpN�N�N�N�N�N�N�N�N OO O0O@OPO`OpO�O�O�O�O�O�O�O�O PP P0P@PPP`PpP�P�P�P�P�P�P�P�P QQ Q0Q@QPQ`QpQ�Q�Q�Q�Q�Q�Q�Q�Q RR R0R@RPR`RpR�R�R�R�R�R�R�R�R SS S0S@SPS`SpS�S�S�S�S�S�S�S�S TT T0T@TPT`TpT�T�T�T�T�T�T�T�T UU U0U@UPU`UpU�U�U�U�U�U�U�U�U VV V0V@VPV`VpV�V�V�V�V�V�V�V�V WW W0W@WPW`WpW�W�W�W�W�W�W�W�W XX X0X@XPX`XpX�X�X�X�X�X�X�X�X YY Y0Y@YPY`YpY�Y�Y�Y�Y�Y�Y�Y�Y ZZ Z0Z@ZPZ`ZpZ�Z�Z�Z�Z�Z�Z�Z�Z [[ [0[@[P[`[p[�[�[�[�[�[�[�[�[ \\ \0\@\P\`\p\�\�\�\�\�\�\�\�\ ]] ]0]@]P]`]p]�]�]�]�]�]�]�]�] ^^ ^0^@^P^`^p^�^�^�^�^�^�^�^�^ __ _0_@_P_`_p_�_�_�_�_�_�_�_�_                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 @@ @0@@@P@`@p@�@�@�@�@�@�@�@�@ AA A0A@APA`ApA�A�A�A�A�A�A�A�A BB B0B@BPB`BpB�B�B�B�B�B�B�B�B CC C0C@CPC`CpC�C�C�C�C�C�C�C�C DD D0D@DPD`DpD�D�D�D�D�D�D�D�D EE E0E@EPE`EpE�E�E�E�E�E�E�E�E FF F0F@FPF`FpF�F�F�F�F�F�F�F�F GG G0G@GPG`GpG�G�G�G�G�G�G�G�G HH H0H@HPH`HpH�H�H�H�H�H�H�H�H II I0I@IPI`IpI�I�I�I�I�I�I�I�I JJ J0J@JPJ`JpJ�J�J�J�J�J�J�J�J KK K0K@KPK`KpK�K�K�K�K�K�K�K�K LL L0L@LPL`LpL�L�L�L�L�L�L�L�L MM M0M@MPM`MpM�M�M�M�M�M�M�M�M NN N0N@NPN`NpN�N�N�N�N�N�N�N�N OO O0O@OPO`OpO�O�O�O�O�O�O�O�O PP P0P@PPP`PpP�P�P�P�P�P�P�P�P QQ Q0Q@QPQ`QpQ�Q�Q�Q�Q�Q�Q�Q�Q RR R0R@RPR`RpR�R�R�R�R�R�R�R�R SS S0S@SPS`SpS�S�S�S�S�S�S�S�S TT T0T@TPT`TpT�T�T�T�T�T�T�T�T UU U0U@UPU`UpU�U�U�U�U�U�U�U�U VV V0V@VPV`VpV�V�V�V�V�V�V�V�V WW W0W@WPW`WpW�W�W�W�W�W�W�W�W XX X0X@XPX`XpX�X�X�X�X�X�X�X�X YY Y0Y@YPY`YpY�Y�Y�Y�Y�Y�Y�Y�Y ZZ Z0Z@ZPZ`ZpZ�Z�Z�Z�Z�Z�Z�Z�Z [[ [0[@[P[`[p[�[�[�[�[�[�[�[�[ \\ \0\@\P\`\p\�\�\�\�\�\�\�\�\ ]] ]0]@]P]`]p]�]�]�]�]�]�]�]�] ^^ ^0^@^P^`^p^�^�^�^�^�^�^�^�^ __ _0_@_P_`_p_�_�_�_�_�_�_�_�_                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                0����������� �����D��   ���� �  XY��x7��� �Ä[��|U�ð��    ����  �����          a2��a2�à��          a2��a2��'��          a2��a2�ç��          a2��a2�ï��           a2��a2�ó��       @   a2��a2�����       �   a2��a2������H���x���            ����     .��   $.��   &.��   9.��   *.��    ..��    1.��   5.��   8.��   ;.��   ?.��   B.��   F.��      @      �H��       ����a2��a2��-X��       \���a2��a2��4X��       ���a2��a2��9X��       ���a2��a2��@X��       t���a2��a2��GX��      ��a2��a2�ûW��      �d��a2��a2��MX��        ��a2��a2�����       <��a2��a2��              h��h��p��p��x��x�À�À�È�È�Ð�Ð�Ø�Ø�à�à�è�è�ð�ð�ø�ø�������������������������������������������������� �� �������������� �� ��(��(��0��0��8��8��@��@��H��H��P��P��X��X��`��`��h��h��p��p��x��x�À�À�È�È�Ð�Ð�Ø�Ø�à�à�è�è�ð�ð�ø�ø�������������������������������������������������� �� �������������� �� ��(��(��0��0��8��8��@��@��H��H��P��P��X��X��`��`��h��h��p��p��x��x�À�À�È�È�Ð�Ð�Ø�Ø�à�à�è�è�ð�ð�ø�ø�������������������������������������������������� �� �������������� �� ��(��(��0��0��8��8��@��@��H��H��P��P��X��X��`��`��h��h��p��p��x��x�À�À�È�È�Ð�Ð�Ø�Ø�à�à�è�è�ð�ð�ø�ø�������������������������������������������������� �� �������������� �� ��(��(��0��0��8��8��@��@��H��H��P��P��X��X��`��`������c��bootargs=root=/dev/mmcblk0p3 rootfstype=ext4 rw console=ttySAC2,115200 bootcmd=movi read kernel 0 40008000;movi read rootfs 0 41000000 100000;bootm 40008000 41000000 bootdelay=3 baudrate=115200 ethaddr=00:40:5c:26:0a:5b ipaddr=192.168.0.20 serverip=192.168.0.10 gatewayip=192.168.0.1 netmask=255.255.255.0   4                                          �e��     �e��   8   �e��      �e��       �e��      �e��      �e��    
  f��    
  gP��      f��	      
f��
              Oj��   Zj��`j��   fj��mj��   h:��tj��   }j�Ãj��   a��G��   �j�Íj��   �j�Ùj������a2��a2��        gi��   ti��zi��   �i�Äi��   �i�Èi��   �i�×i��   �i�ái��   �i�ñi��   �i���i��   �i���i��   �i���i��   �i���i��   �i���i��   �i�� j��	   �Y��	j��
   j��j��   j��$j��   1j��:j��   Cj��Ij������a2��a2��        �h��   p�Ôh��   �h�îh��   v�÷h��   �h���h��   '���h��   	���h��   �h���h��   i��i��	   'i��0i��
   Di��Mi������a2��a2��    �I��%h��   2h��8h��   Ih��Nh��   ^h��ch��   sh��wh������a2��a2��              �����S�èS�ïS������'  �� @B ���     
                     #   (   -   2   7   <   F   P   s5pser0         S5PUART0����    ����������������$���    s5pser1         S5PUART1���    ����������������    s5pser2         S5PUART2$���    ,���4���<����������    s5pser3         S5PUART3D���    L���T���\��ü������             �����������������������������������~������~          bootloader                             recovery                 P             kernel            `       P             ramdisk           �       0             system            �       �           cache             �                  userdata          �                         ��������   ����/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               (((((�AAAAAABBBBBB                                �����������  �����  �  
   
      �              u��      �d��|��a2�����       f�������g��       �d��m��a2��;��      �q��A��d��c��      h��m��a2�Ï��      h��m��a2�Õ��      �g�Ü��������      �u�������1��      4u��8��U�ÿ��      v�����a2��Z0��      w���������       H{����@�é��       |x�ð��������      �|����a2�ü��      4���������J��       �}��S��{����       �}��"��D�Û��       �}�æ�����"(��      ����+(��P(��b+��       ����j+�Ü+��8,��      ����������>,��      ����F,��s,���,��       ̢���,���,��Q-��      H���V-��v-���-��      H����-��a2��I.��       ����O.��t.�á0��       ��ç0���0��1��       ȯ��1��E1���.��       ȯ�ä1��E1��S��      (��â3�ñ3���3��      ����3��4��4��      ���4��4��;4��      ���>4��R4��u4��      ����x4�Ä4�å4��      P��é4�ø4���4��      �����4���4��35��      ����85��T5���5��      �����5���5��6��      ���6��/6��T6��       ���Z6��x6�Ù:��       ���á:��a2���:��       \����:���:���:��      T���i;��x;��>��       ����>��8>��	@��       l���@��:@�ÿJ��       ����J���J���F��       ����K��:K�ÛP��      ���áP���P���P��      ����Q���P��0Q��      ����4Q���P��^Q��      @���cQ�ÊQ�ÂT��        �ÊT��a2�ÆT��      ���ûT���T��AV��       ���IV��cV�ÏV��      �ØV�ôV�ù&��       <��(W��BW�ûW��      �d�ÿW���W��RX��      ��ZX��a2��
Y��       P	��Y��(Y��*6��      �	�ÂY�ÜY�åY��      �	�ëY��    �Y��      �	���Y��    �]��      p�ï]�þ]��Z^��       P��^^�ò^�ö���      `���^��a2���_��      ����_��`��Ne��      �>��Ve��ve��  ��   $ ��   ( ��   , ��   0 ��   4 ��   8 ��   ���   ���   	��   ���   ��   8��   <��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��    ��   �$��   �$��    %��   l'��   �'��   �'��   �'��   �'��   (��   <(��   X(��   �(��   �(��   �(��   �(��   $)��   P)��   l)��   �)��   �)��   �)��   *��   $*��   L*��   �*��   �*��   �*��   �*��   +��   D+��   x+��   �+��   �+��   �+��   ,��   <,��   p,��   �,��   �,��   �,��   -��   4-��   h-��   �-��   �-��   �-��   .��   ,.��   `.��   �.��   �.��   �.��   �.��   $/��   X/��   x/��   �/��   �/��   �/��   0��   P0��   p0��   �0��   �0��   �0��   1��   H1��   d1��   �1��   �1��   �1��   �1��   2��   ,2��   L2��   t2��   �2��   �2��   �2��   �2��   3��   <3��   X3��   x3��   �3��   �3��   �3��   4��    4��   @4��   h4��   �4��   �4��   �4��   �4��   5��   05��   L5��   l5��   �5��   �5��   �5��   �5��   6��   46��   \6��   �6��   �6��   �6��   7��   7��   47��   L7��   d7��   �7��   �7��   �7��   �7��   ,8��   48��   d8��   L9��   P9��   T9��   P:��   T:��   X:��   X;��   \;��   `;��   @<��   D<��   H<��   (=��   ,=��   0=��   �=��   �=��   �=��   �>��   �>��   �>��   �?��   �?��   �?��   �@��   �@��   �@��   �A��   �A��   �A��   �B��   �B��   �B��   �C��   �C��   �C��   �D��   �D��   �D��   �E��   �E��   �E��   �F��   �F��   �F��   �G��   �G��   �G��   �H��   �H��   �H��   �I��   �I��   �I��   |J��   �J��   �J��   hK��   lK��   pK��   TL��   XL��   \L��   @M��   DM��   HM��   ,N��   0N��   4N��   �N��   �N��   �N��   �O��   �O��   �O��   �P��   �P��   �P��   �Q��   �Q��   �Q��   �R��   �R��   �R��   pS��   tS��   xS��   DU��   HU��   LU��   PU��   TU��   XU��   \U��   `U��   dU��   hU��   xU��   �U��   �U��   �W��   �Y��   �Y��   Z��   lZ��    [��   �[��   �[��   �[��   �\��    ]��   ]��   ]��   ]��   ]��    ]��   $]��   (]��   �]��   �]��    ^��   ^��   ^��   ^��   ^��   ^��    `��   $`��   (`��   ,`��   4`��   <`��   H`��   b��   Dc��   Hc��   Lc��   Pc��   Tc��   Xc��   \c��   `c��   dc��   hc��   �c��   �c��   �c��   �c��   d��   8d��   \d��   �d��   �d��   �d��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��   �e��    f��   f��   �f��   �f��   �g��   �g��   �g��   �g��   �g��   �g��   �g��   �g��    h��   0h��   hh��   �h��   i��   hi��   li��   �j��   �j��   �j��   �j��   �j��   �j��   �j��   �k��   �k��   �k��   <o��   @o��   Do��   Ho��   Lo��   Po��   To��   Xo��   \o��   `o��   do��   ho��   lo��   po��   to��   xo��   |o��   �q��   �q��   �q��   �q��   �q��   �q��   �q��   �q��   �q��   �q��   �t��   �t��   �t��   �t��   �t��   �t��   �t��   �t��   �t��   �t��   �t��   ,u��   0u��   �u��   �u��   �u��   v��   v��   v��   �v��   �v��    w��   w��   w��   �w��   �w��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��   �z��    {��   �|��   �|��   �|��   �}��   �}��   �}��   �}��   �}��   �}��   �}��   ~��   ~��   ~��   ~��   ���   ����   ���   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   P���   T���   X���   \���   `���   d���   ����   ����   Ă��   8���   h���   l���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ���   ܉��   ����   ���   ���   ���   ����   ���   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   \���   `���   d���   h���   l���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ĕ��   ȕ��   ̕��   Е��   ԕ��   ؕ��   ܕ��   ����   ���   ���   ���   ���   ����   ����   ����    ���   <���   @���   D���   ����   ����   ����   ����   ġ��   ȡ��   ̡��   С��   ԡ��   ء��   ܡ��   ���   ���   ���   ���   ���   ����   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   H���   L���   P���   T���   X���   \���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   Ģ��   Ȣ��   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   $���   (���   ,���   0���   4���   8���   <���   @���   D���   ����   ����   ����   Ĩ��   Ȩ��   ̨��   Ш��   Ԩ��   L���   P���   T���   X���   \���   `���   ���   ����   ����   4���   8���   <���   @���   D���   H���   L���   ����   ���   ���   0���   P���   l���   ����   ���   ܭ��   8���   <���   ����   ����   ����   ����   ����   ����   ����   ���   ����   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ���   ���   ���   ���   ���   ���   ���   ���   ���   ����   ����   ����   ����   ܷ��   ���   p���   t���   x���   |���   ����   H���   L���   ����   ����   ļ��   ȼ��   ̼��   м��   Լ��   ؼ��   ܼ��   ���   ����   ̾��   о��   Ծ��   ؾ��   ܾ��   ���   ���   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   H���   L���   P���   l���   p���   t���   x���   |���   ����   ����   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   H���   L���   P���   T���   X���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   x���   |���   ����   ����    ���   ���   ����   ����   ����   ����    ���   ���   ����   \���   `���   d���   h���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   ���   ���   ����   H���   L���   P���   T���   ����    ���   ���   ���   X���   \���   `���   d���    ���   ���   ���   ���   ���   ���   4���   8���   ����   <���   @���   D���   H���   L���   P���   ����   ����   ����   ����   ����   ����   ����    ���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   X���   \���   `���   d���   h���   l���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ���   @���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   ���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   ����   ����   ����   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   X���   p���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ��   4 ��   8 ��   ��   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   0	��   4	��   <	��   @	��   D	��   H	��   L	��   �	��   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   T��   X��   \��   `��   d��   h��   l��   p��   t��   x��   ��   ��   ��   ��    ��   $��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   P��   T��   X��   \��   `��   d��   h��   ���    ��   $��   (��   ,��   0��   ���   ���   ���   ���   ���   ���   ���   ���   l��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   @��   D��   H��   L��   P��   T��   x��   |��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   P��   T��   X��   ���   ���    ��   ��   ���   ���   H��   L��   ���   ���    ��   < ��   h ��   � ��   � ��   � ��   � ��   �"��   �"��   �"��   �"��   �"��   �"��   �"��   �"��   �#��   �#��   �$��   �%��   �%��   �%��   �%��   �%��   �%��   l&��   p&��   t&��   �&��   �&��   �&��   �&��   $'��   ('��   X'��   �'��   |(��   �(��   �*��   �*��   �*��   �0��   �0��   �0��   �0��   �2��   h7��   �7��   8��   8��   8��    8��   $8��   x8��   �8��   P9��   T9��   X9��   �9��   �9��   `:��   d:��   h:��   l:��   p:��   t:��   x:��   �:��   X;��   \;��   `;��   d;��   h;��   l;��   �;��   ,=��   0=��   4=��   8=��   <=��   @=��   D=��   H=��   L=��   P=��   T=��   X=��   \=��   `=��   d=��   h=��   l=��   p=��   �=��   @>��   D>��   T>��   �>��   �>��   �>��   �?��   �?��   �?��   �?��   @��   @��    @��   @@��    B��   $B��   (B��   ,B��   0B��   �C��   �C��   �C��   4F��   8F��   TI��   XI��    K��   K��   K��   K��   lK��   pK��   tK��   xK��   |K��   @L��   �Q��    R��   R��   R��   R��   R��   PR��   TR��   S��   �Z��   �Z��   �Z��    [��   [��   [��   �[��   �[��   �[��   �[��   �[��   �[��   �[��   �[��   T\��   �\��   �\��   �\��   �\��   �\��   �\��   �\��    ]��   �]��    ^��   p_��   t_��   x_��   |_��   �_��   �_��   �_��   �_��   �_��   �_��   �`��   �`��   �`��   �`��   $a��   (a��   �c��   �c��   �c��    d��   d��   d��   d��   d��   d��   d��   �d��   e��   �h��   �h��   �h��   �h��   �i��   �i��   �j��   xl��   |l��   �l��   �l��   �l��   �l��   �l��   �l��   ,s��   0s��   4s��   8s��   <s��   @s��   Ds��   Hs��   Ls��   hs��   Pt��   Tt��   Xt��   \t��   Dv��   Hv��   Lv��   Pv��   Tv��   Xv��   \v��   `v��   dv��   hv��   Hx��   hx��   �x��   �x��   y��   Ty��   �y��   �y��   $z��   pz��   �z��   �z��   �z��   �z��   <{��   H{��   �{��   �{��   $|��   �|��   �|��   �|��   �|��   �|��   �|��   �|��   �}��   ~��   D~��   H~��   �~��   �~��   �~��   4���   p���   t���   ā��   ȁ��   ́��   d���   ���   P���   T���   ،��   ܑ��   ����   ���   ���   ���   ���   X���   \���   `���   d���   В��   Ԓ��   ؒ��   ܒ��   ����   8���   <���   ����   ����   ����   ����   ���   ���   P���   X���   \���   `���   d���   ����   P���   T���   X���   ���   <���   @���   D���   H���   L���   P���   T���   X���   ĝ��   ȝ��   ̝��   Н��   ԝ��   ؝��   ܝ��   ����   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   ���   ���   ���   ����   ����   ����    ���   ���   ğ��   ȟ��   ̟��   П��   ԟ��   ؟��   ܟ��   ����   ���   ���   ���   ���   ����   ����   ����    ���   ���   ����   ����   ����   ����   ����   ����   ����   ����   ܢ��   ���   ���   ���   ���   ���   ����   ����   ���   ���   ���   ���   ����   ����   ����    ���   ,���   ����   ����   ����   Į��   Ȯ��   ̮��   Ю��   Ԯ��   خ��   ܮ��   ���   ���   H���   L���   P���   T���   ����   ����   ���   ���   ���   ����   ����   ����    ���   ���   ����   ����   ����   İ��   Ȱ��   ̰��   а��   ԰��   ذ��   ����   ����   ����   ����   ����   Ĳ��   Ȳ��   ̲��   в��   Բ��   ز��   ܲ��   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ����   ����   ����   ����   ����   d���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   D���   H���   L���   P���   ����   ����   ����   ����   ����    ���   ���   ����   ����   ����   ����   ����   ����   ���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   ���   ����   ����   ����   ����   ����   ����   ����   ����   H���   p���   t���   ����   ����   (���   ,���   0���   ����   ����   ����   (���   d���   ����   (���   ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   ���   ���    ���   ���   ���   ���   ���   ���   ����   ����   ���   0���   8���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ���    ���   |���   ����   x���   ���   ���   ���   ���    ���   $���   (���   x���   |���   ����   ����   ���   ����   ���   ����   ����   (���   x���   ����   ����   ����   ���   l���    ���   ���   ���   ���   ���   ���   X���   \���   `���   ����   ���   ���   ���   ���   ���    ���   $���   ����   ����   ����   ����   X���   `���   ����   p���   ����   L���   ����   ����   l���   p���   ����   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   8���   ����   ����   ����   ����    ���   ����   ����   ����   ����   ����   ����   ����   ����   0 ��   � ��   P��   T��   X��   \��   `��   d��   ���   ��   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   P��   T��   X��   \��   `��   d��   h��   l��   d-��   h-��   l-��   p-��   �-��   @.��   D.��   �/��   �/��   x4��   |4��   �4��   �4��   �4��   �4��   �4��   �4��   �4��   �4��   47��   87��   <7��   @7��   D7��   �9��   H:��   �:��   L;��   P;��   =��   =��   =��    =��   $=��   (=��   t=��   �=��   �A��   �A��   �A��    B��   B��   B��   B��   B��   B��   �B��   �B��   �B��   �B��   �B��   �B��   �B��   �B��   �B��   �B��    C��   C��   C��   C��   `E��   dE��   \O��   `O��   dO��   hO��   lO��   pO��   tO��   �O��   �O��   �O��   �O��   �O��   �P��   �P��   �P��    Q��   Q��   Q��   Q��   �V��   �V��   �V��   �V��   �V��   �V��   �V��   �V��   �V��   �V��   �V��   �V��    W��   W��   W��   W��   W��   W��   W��   W��    W��   $W��   (W��   ,W��   0W��   4W��   8W��   <W��   @W��   DW��   HW��   LW��   dW��   �W��   �W��    X��   X��   �X��   �X��   �X��   �X��   �X��   �X��   �X��   �Z��   �Z��   �Z��   �Z��   ([��   \��   ]��   ]��   ]��   ]��   4]��   8]��   �^��   �^��   �^��   �^��   t`��   x`��   |`��   �`��   �`��   4a��   8a��   �a��   �a��   xb��   �b��   �d��   �d��   �d��   �g��   @h��   Lh��   �j��   �j��   �j��   �j��   tp��   Tu��   �x��   �x��   y��   8y��   �y��   p{��   `}��   ����   ����   ����   ����   ����    ���   d���   h���   ����   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   H���   L���   P���   T���   X���   \���   `���   d���   h���   l���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   8���   <���   @���   D���   H���   L���   P���   ���   ���   ���   ���    ���   $���   (���   0���   4���   8���   <���   @���   D���   H���   L���   P���   T���   X���   \���   `���   d���   d���   h���   l���   p���   t���   x���   |���   ����   ����   ����   ĳ��    ���   d���   ����   ���   ���   D���   `���   d���   ����   X���   \���   ����    ���   ���   ���   ���   ����   ����   Է��   ����   ����   P���   T���   Ļ��   Ȼ��   ̻��   л��   Ի��   ػ��   ܻ��   ���   ���   ���   ���   ���   ����   ����   ����    ���   ���   ���   ���   ���   4���   H���   ����   ܽ��   ���   (���   t���   `���   ���   ���   P���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ���   D���   H���   d���   T���   X���   \���   `���   d���   h���   l���   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   p���   t���   x���   |���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   4���   ����   |���   ����   ����   ����   ����   ����   ����   ����   ���   h���   ����   ����   ����   ����   ����   ����   ����   ����    ���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ���   ���   @���   D���   L���   P���   T���   ����   ����   ����   ����   ����   ����   ����   ���   ���    ���   $���   (���   ,���   0���   4���   8���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   `���   d���   h���   l���   p���    ���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ,���   0���   4���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����    ���   ���   ���   ���   ���   ���   (���   L���   T���   \���   l���   ���   ���   ���   ���   ���   ���   ���    ���   $���   (���   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ����   ,���   0���   4���   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   ( ��   , ��   0 ��   4 ��   8 ��   < ��   L ��   \ ��   ` ��   d ��   t ��   x ��   | ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   � ��   ��   ��   $��   ,��   4��   <��   D��   L��   T��   \��   d��   l��   t��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   $��   (��   ,��   0��   <��   @��   D��   H��   T��   X��   \��   p��   t��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   P��   T��   X��   \��   `��   d��   h��   l��   p��   t��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   P��   T��   X��   \��   `��   d��   h��   l��   p��   t��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   P��   T��   X��   \��   `��   d��   h��   l��   p��   t��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   ��   ��    ��   $��   (��   ,��   0��   4��   8��   <��   @��   D��   H��   L��   P��   T��   X��   \��   `��   d��   h��   l��   t��   ���   ���   ���   ���   ��   ��    ��   ,��   8��   D��   P��   d��   l��   p��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    	��   	��   	��   	��   	��    	��   $	��   ,	��   0	��   8	��   <	��   D	��   H	��   P	��   T	��   \	��   `	��   h	��   l	��   t	��   x	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   �	��   
��   
��   
��   
��   
��    
��   (
��   ,
��   4
��   8
��   @
��   D
��   L
��   P
��   X
��   \
��   d
��   h
��   p
��   t
��   |
��   �
��   �
��   �
��   �
��   ��   ��   ��    ��   $��   (��   H��   P��   T��   X��   \��   `��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��    ��   $��   0��   4��   8��   <��   H��   L��   P��   T��   `��   d��   h��   l��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��   ��   ��   ��    ��   $��   (��   ,��   8��   <��   @��   D��   P��   T��   X��   \��   h��   l��   p��   t��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   (��   ,��   0��   4��   @��   D��   H��   L��   X��   \��   `��   d��   p��   t��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��    ��   $��   0��   4��   8��   <��   H��   L��   P��   T��   `��   d��   h��   l��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��   ��   ��   ��    ��   $��   (��   ,��   8��   <��   @��   D��   P��   T��   X��   \��   h��   l��   p��   t��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���    ��   ��   ��   ��   ��   ��   (��   ,��   4��   @��   D��   L��   X��   \��   `��   d��   p��   t��   x��   |��   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���                         ��            ��      %   ���     	    |��     ��   ���     ��R   ���      C   4{��     
     �=��      5   4{��     	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ������  ���������������������D   �����!� P�  
 P�  
  P�   
����O�@�  �џ� -�r  ���0�  �џ��  �  P��M @��� -���0�  �tџ� -�� �   �  �`џ��  �  P��M @��� -�  �A  �� ��% ��� @�@��@�� ���o���?P�T���� ��0�Q�0/�?�0O�? ��?��?P�$���� ��? ��0�Q�0/�?�0O�?��                                                                                                                                 ���0 ��0�� ���� ���� ���O��o���� � � ��?   � � � ��-� ����M� ��2�� 0��� �1 �2@�  ��0� 0��S�  0�P ��S<�S9D� R�   
����0�@ ��(0 �2@�  ��0�D ��(0 �2@� ��0�H ��(0 �2@� ��0�L ��(0 �2@� �� 0 �2@�   �p A�  �� 0 �2@�(�� �� 0 �2@� �� �� 0 �2@� �� �� 0 �2@�   � A� �� 0 �2@�(�� �� 0 �2@� �� �� 0 �2@�   �H A� �� 0 �2@�   �I A�  �� 0 �2@� ��$ �� 0�� �� Ћ� ���/�e p�  
 p�l  
 p�k  
 p�n  
 p�  
 p�  
 p�  
 p�  
 p�  
 p�  
 p�  
 p�  
�  �P�  
P�8  
��� P�0/�  
�� P�/�  
��� P�0/�  
���� P�  ��  
��� P�  ��  
��� P�  ��  
��� P�  ��  
��� P�  ��  
x�� P�  ��  
l�� P�  ��  
`�� P�  ��  
T�� P�  ��  
H�� P�  ��  
<�� P�  �~  
���� P�  �y  
��� P�  �u  
��� P�  �q  
��� P�  �m  
��� P�  �i  
��� P�  �e  
b  �d  �  ���� ��0��_  ��_-����� ����� �� ������ �� ������  �� ��  ���� ��  �� ��  ������$X��P�,���  �  P�  O��� �X��(X���_��  �� ��  �� 0��8  �<�����4�� �� ��� �/  � @-���� @������!��  ��  ��!��  ��  ��O��� �!  ��0/�  �� �� ��  �� ����!��`?��  �� �����������  � ����|��|7�� �  R���� ��0��  � ��@��  �����  ����  ����  <  @/P0 `0 a4 `4 a !P!P!P`/P�/P!P ` a �� 	�  `�    4$   4 �  P��  �-� ����M� �� �4 �0A�  ��  �� 4 �0A� ��  ��$4 �0A�  ��  ��(4 �0A�  ��  ��,4 �0A�  ��  ��0��0� 4 �0A� �  ��4 �0A� 0��0�0�0�  S�   0��Z  �04 �0A�   � A�  ��  ��44 �0A�  � A�  ��  ��84 �0A�  � A�  ��  ��<4 �0A�  � A�  ��  ��@4 �0A� �  ��4 �0A� 0��0�0�@0�  S����
4 �0A�@ ��  ��0�0� 5 �0A�  ��0�  ��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0�0�5 �0A�  ��0�  ��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0�� 0�� �� Ћ� ���/� H-����8�M� 0�2@�0�(0 �2@�0��0�(0 �2@�0��':��0�':��0�( K�80K� ����  ��/O�^��� 0��  S�  
 0��9 �2 �0A� 0��0�0�0�  S�  
 0��/ �4 �0A� 0��0�0�0�  S�   0��% �(0 �0A� ��  ��80 �0A� ��  ��0 �0A� ��  ��0��0�0�0��0�0�
=��0�0�;��0� 2 �0A� �  ��0��0�0�0��0�4 �0A� �  ��2 �0A�( �  ��2 �0A�$ �  ��2 �0A�  �  ��2 �0A� �  ��02 �0A�8 �  ��42 �0A�4 �  ��82 �0A�0 �  ��<2 �0A�, �  ��p4 �0A�( �  ��t4 �0A�$ �  ��x4 �0A�  �  ��|4 �0A� �  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A�  ��  ��4 �0A� ��  �� 4 �0A� �  ��$4 �0A�  ��  ��(4 �0A�  ��  ��,4 �0A�  ��  ��0��0� 4 �0A� �  ��00 �0A� �  ��40 �0A� �  �� 0 �0A� �  ��$0 �0A� �  ��0 �0A� 0��0�0�0�  S����
0 �0A� ��  ��2 �0A�  ��  ��2 �0A�  ��  ��2 �0A�  ��  ��2 �0A�  ��  ��02 �0A�  ��  ��42 �0A�  ��  ��82 �0A�  ��  ��<2 �0A�  ��  ��4 �0A� 0��0�0�@0�  S����
4 �0A�@ ��  ��p4 �0A�  ��  ��t4 �0A�  ��  ��x4 �0A�  ��  ��|4 �0A�  ��  �� 5 �0A�  ��0�  ��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0��0� ��5 �0A� 0�� 0�� 0�� ���K� ����-� ����M� � 0 �2@� 0��0� 0��0�0�0��  ��0�  ��0�0��  ��0� ��0�0��  ��0� ��0�00��  ��0� ��0�40��  ��0� �� 0��0�/  �0� �"���� � ��,��  ��� ��0�� ����0��  ��0� �"���� � ��A/��  ��� ��0�� ����0��  ��0� �"���� � ��B/��  ��� ��0�� ����0��  ��0�0��0� � 0 �2@�0�� R����: 0�� �� Ћ� ���/��-� ����M� � 0 �2@� 0��0� 0 �2@�0��0� 0��0� 0��0� 0��0�X  �0�0�� �  ��  ��0�0�� � ��  ��0�0�� � ��  ��0�00�� � ��  ��0�40�� � ��  �� 0��0�/  �0�2�� ��0�0��<�� �� �� �� ���� ��  ��  ��0�2�� ��0�0��A?�� �� �� �� ���� ��  ��  ��0�2�� ��0�0��B?�� �� �� �� ���� ��  ��  ��0�0��0� � 0 �2@�0�� R����: �0�0��0�0�0��0� � 0 �2@�0�� R���: 0�� �� Ћ� ���/��-� ����M� � 0 �2@�0��0� 0 �2@�0��0� 0��0�0�  ��0�  �� 0��0�5  � �0�;��  ���0�� ����0��  �� �0�;��0��  ���0�� ����0��  �� �0�>��0��  ���0�� ��0������0��  �� �0�>��0��  ���0�� ��0������0��  �� �0�0��0�0�0��0� � 0 �2@�0�� R����: 0�� �� Ћ� ���/��-� ����M� � 0 �2@�0��0� 0 �2@�0��0� 0��0�0� �  ��  �� 0��0�H  �0�;��0��  ��  ��0�;��0�� �� �� ���� ��  ��  ��0�>��0��  ��  ��0�>�� �� �� ���� ��  ��  ��0�>��  ��  ��0�>��0�� �� �� �� ������ ��  ��  ��0�>��0��  ��  ��0�>��0�� �� �� �� ������ ��  ��  �� �0�0��0�0�0��0� � 0 �2@�0�� R���: 0�� �� Ћ� ���/��-� ����M� � 0 �2@�0��0� 0 �2@� 0��0� 0 �2@�$0��0��2��0� 0��0�0�  ��0�  ��0�0��  ��0� ��0�0��  ��0� ��0�  ��0� �� 0��0�  � �0�1����0�0���0�� ��0� ����0�0��0� �0� R����� 0��0�  � �0�1����0�0��<�� ��0� ����0�0��0� �0� R����� 0�� �� Ћ� ���/��-� ����M� � 0 �2@�0��0� 0 �2@� 0��0� 0 �2@�$0��0��2��0� 0��0�0� �  ��  ��0�0�� � ��  ��0�0�� � ��  ��0� � ��  �� 0��0�  �0�1�� ��0�0���0��� ���!��  ��0�0��0� �0� R����� 0��0�  �0�1�� ��0�0��=��  ��  ��0�1�� ��0�0��<��� ����� � � �� !�� �� �  ��0�0��0� �0� R����� 0�� �� Ћ� ���/� H-����8  �@���� ����� ��>��� 0�� �� ���| @ H-�����M� �8  �@����� ������ ����� 0�� ���K� ���| @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                !1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������!1AQaq��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                @@!@1@A@Q@a@q@�@�@�@�@�@�@�@�@AA!A1AAAQAaAqA�A�A�A�A�A�A�A�ABB!B1BABQBaBqB�B�B�B�B�B�B�B�BCC!C1CACQCaCqC�C�C�C�C�C�C�C�CDD!D1DADQDaDqD�D�D�D�D�D�D�D�DEE!E1EAEQEaEqE�E�E�E�E�E�E�E�EFF!F1FAFQFaFqF�F�F�F�F�F�F�F�FGG!G1GAGQGaGqG�G�G�G�G�G�G�G�GHH!H1HAHQHaHqH�H�H�H�H�H�H�H�HII!I1IAIQIaIqI�I�I�I�I�I�I�I�IJJ!J1JAJQJaJqJ�J�J�J�J�J�J�J�JKK!K1KAKQKaKqK�K�K�K�K�K�K�K�KLL!L1LALQLaLqL�L�L�L�L�L�L�L�LMM!M1MAMQMaMqM�M�M�M�M�M�M�M�MNN!N1NANQNaNqN�N�N�N�N�N�N�N�NOO!O1OAOQOaOqO�O�O�O�O�O�O�O�OPP!P1PAPQPaPqP�P�P�P�P�P�P�P�PQQ!Q1QAQQQaQqQ�Q�Q�Q�Q�Q�Q�Q�QRR!R1RARQRaRqR�R�R�R�R�R�R�R�RSS!S1SASQSaSqS�S�S�S�S�S�S�S�STT!T1TATQTaTqT�T�T�T�T�T�T�T�TUU!U1UAUQUaUqU�U�U�U�U�U�U�U�UVV!V1VAVQVaVqV�V�V�V�V�V�V�V�VWW!W1WAWQWaWqW�W�W�W�W�W�W�W�WXX!X1XAXQXaXqX�X�X�X�X�X�X�X�XYY!Y1YAYQYaYqY�Y�Y�Y�Y�Y�Y�Y�YZZ!Z1ZAZQZaZqZ�Z�Z�Z�Z�Z�Z�Z�Z[[![1[A[Q[a[q[�[�[�[�[�[�[�[�[\\!\1\A\Q\a\q\�\�\�\�\�\�\�\�\]]!]1]A]Q]a]q]�]�]�]�]�]�]�]�]^^!^1^A^Q^a^q^�^�^�^�^�^�^�^�^__!_1_A_Q_a_q_�_�_�_�_�_�_�_�_``!`1`A`Q`a`q`�`�`�`�`�`�`�`�`aa!a1aAaQaaaqa�a�a�a�a�a�a�a�abb!b1bAbQbabqb�b�b�b�b�b�b�b�bcc!c1cAcQcacqc�c�c�c�c�c�c�c�cdd!d1dAdQdadqd�d�d�d�d�d�d�d�dee!e1eAeQeaeqe�e�e�e�e�e�e�e�eff!f1fAfQfafqf�f�f�f�f�f�f�f�fgg!g1gAgQgagqg�g�g�g�g�g�g�g�ghh!h1hAhQhahqh�h�h�h�h�h�h�h�hii!i1iAiQiaiqi�i�i�i�i�i�i�i�ijj!j1jAjQjajqj�j�j�j�j�j�j�j�jkk!k1kAkQkakqk�k�k�k�k�k�k�k�kll!l1lAlQlalql�l�l�l�l�l�l�l�lmm!m1mAmQmamqm�m�m�m�m�m�m�m�mnn!n1nAnQnanqn�n�n�n�n�n�n�n�noo!o1oAoQoaoqo�o�o�o�o�o�o�o�opp!p1pApQpapqp�p�p�p�p�p�p�p�pqq!q1qAqQqaqqq�q�q�q�q�q�q�q�qrr!r1rArQrarqr�r�r�r�r�r�r�r�rss!s1sAsQsasqs�s�s�s�s�s�s�s�stt!t1tAtQtatqt�t�t�t�t�t�t�t�tuu!u1uAuQuauqu�u�u�u�u�u�u�u�uvv!v1vAvQvavqv�v�v�v�v�v�v�v�vww!w1wAwQwawqw�w�w�w�w�w�w�w�wxx!x1xAxQxaxqx�x�x�x�x�x�x�x�xyy!y1yAyQyayqy�y�y�y�y�y�y�y�yzz!z1zAzQzazqz�z�z�z�z�z�z�z�z{{!{1{A{Q{a{q{�{�{�{�{�{�{�{�{||!|1|A|Q|a|q|�|�|�|�|�|�|�|�|}}!}1}A}Q}a}q}�}�}�}�}�}�}�}�}~~!~1~A~Q~a~q~�~�~�~�~�~�~�~�~!1AQaq����������!�1�A�Q�a�q�����������р����!�1�A�Q�a�q�����������с����!�1�A�Q�a�q�����������т����!�1�A�Q�a�q�����������у����!�1�A�Q�a�q�����������ф����!�1�A�Q�a�q�����������х����!�1�A�Q�a�q�����������ц����!�1�A�Q�a�q�����������ч����!�1�A�Q�a�q�����������ш����!�1�A�Q�a�q�����������щ����!�1�A�Q�a�q�����������ъ����!�1�A�Q�a�q�����������ы����!�1�A�Q�a�q�����������ь����!�1�A�Q�a�q�����������э����!�1�A�Q�a�q�����������ю����!�1�A�Q�a�q�����������я����!�1�A�Q�a�q�����������ѐ����!�1�A�Q�a�q�����������ё����!�1�A�Q�a�q�����������ђ����!�1�A�Q�a�q�����������ѓ����!�1�A�Q�a�q�����������є����!�1�A�Q�a�q�����������ѕ����!�1�A�Q�a�q�����������і����!�1�A�Q�a�q�����������ї����!�1�A�Q�a�q�����������ј����!�1�A�Q�a�q�����������љ����!�1�A�Q�a�q�����������њ����!�1�A�Q�a�q�����������ћ����!�1�A�Q�a�q�����������ќ����!�1�A�Q�a�q�����������ѝ����!�1�A�Q�a�q�����������ў����!�1�A�Q�a�q�����������џ����!�1�A�Q�a�q�����������Ѡ����!�1�A�Q�a�q�����������ѡ����!�1�A�Q�a�q�����������Ѣ����!�1�A�Q�a�q�����������ѣ����!�1�A�Q�a�q�����������Ѥ����!�1�A�Q�a�q�����������ѥ����!�1�A�Q�a�q�����������Ѧ����!�1�A�Q�a�q�����������ѧ����!�1�A�Q�a�q�����������Ѩ����!�1�A�Q�a�q�����������ѩ����!�1�A�Q�a�q�����������Ѫ����!�1�A�Q�a�q�����������ѫ����!�1�A�Q�a�q�����������Ѭ����!�1�A�Q�a�q�����������ѭ����!�1�A�Q�a�q�����������Ѯ����!�1�A�Q�a�q�����������ѯ����!�1�A�Q�a�q�����������Ѱ����!�1�A�Q�a�q�����������ѱ����!�1�A�Q�a�q�����������Ѳ����!�1�A�Q�a�q�����������ѳ����!�1�A�Q�a�q�����������Ѵ����!�1�A�Q�a�q�����������ѵ����!�1�A�Q�a�q�����������Ѷ����!�1�A�Q�a�q�����������ѷ����!�1�A�Q�a�q�����������Ѹ����!�1�A�Q�a�q�����������ѹ����!�1�A�Q�a�q�����������Ѻ����!�1�A�Q�a�q�����������ѻ����!�1�A�Q�a�q�����������Ѽ����!�1�A�Q�a�q�����������ѽ����!�1�A�Q�a�q�����������Ѿ����!�1�A�Q�a�q�����������ѿ����!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�������������������!�1�A�Q�a�q�����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                